��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������r��#@�/�����4�p5���4;Od��N��r�I#��7h��$�(��?�g:�ZGY�bӍ��0Yzb0o �Β��A���p�6� �����4���e��Ǟ�H� �a�C���t.����+^���}��G�|lm�.�|����"��(�cx�m1�#�N�N�:k?n~Sn`�'|���y1/)�
x@���n�+J�\O{&	�.�B䛄�%��i�f�f�L�u��i/���R�@;C�!�M*.ɪ ��_�zG�ȍ��ڸA�9[Íp���="N�jZ��|݈��y�A���_�������ⳤ\B�ҥL������x%��}�D��c��t�s����PF`�t|����Nl��W�`f2�C3�$�IF��<�Χ�[���jY9 �$Rv3�4H�6\�&�;��n�7WJ�Q(��KB���"V�� �z���0S��:�A�m�M�WX4�ip5(p���q���r�y|��[��cᰙ"�G�_:-����$IE-2����Tg$�����!�M��A ��
Xm�b}O !�N�w:QP�!��7+1�G�*FzL}��sce�'�ы��[_��4�'׆P�����5�J/A@�>�+<����g|(�Aem[z(���%���2I'�:�S�vHv�wL��U W�!��qѾ�+��9����-+�l:��6?f>�9i�ԕ�l>ʛ���e������8&�ԟ.6��x�n�C_򧊎�&��c"�#`���O|��$M;&�Ā(%����>l����೧+���cp"�%�L�[�Bs�-o�0)I�O�:���tea��hÿ�j�)/�C���nK���8��֚UH���(�C�#�������)��I�2ڵ7���V���
%2 \� {��Dv��ݲ�1�<�_X������{�,�����L?�/��3=�!�4���]RRo�l�IV�E���7%�l�
��+c����B��3�2|,U�A�����̷��3l�PK8�Od#���ǋM�����`��������g~V=��X�x�vVӑ,$� ����Qb���zj����͆�0t�R(�y�'3@���H:NW����g"�z��/ ����?�����C�en�]�������,�͹u^C�� �<��$��h"��!��d��� !X5r?�ޥG�����ʉ����֨͛�2@��o0� [be��-�r�e�M�E��rӀ�=M+��yN^�P���@���N(M��>�#me�GorX��&1�8+_�3�gx�Z	�#��oy��X�v/�Gg�V[/#����R��c+g�1�s6�Y�EL�C�g��)8�۰G1��A�'i��s�Q�W�od])���7��e����)�;;���*���h�ׯ�_��[Q�.ƈ�Q0�4���'i���]�FO�z��;�D>�%�>΢����D�+x�%���s����N��m���!�ͥ�e�ŏ�O%E�Zj_��0�E���=L�V�	|��P]`&�T�|Ɖ�g+����E�}�Q����U0����y0Ǧo��"حt9�&���V0�9�;��1�D�婠iGT�6܂Io$�RR� ��ͪ�U���4��Do/�l&����'�
즚��[q5@�0���8�D;��Ht�%�^֥�F۠���|3R���gEh������H?Q��N�ic_S6f�����_�M�͸�Vɉ��M�s��h�|;��K���^��ġD�\����֚����Mt<pBO<)%3@�g/9�F��i�.��jCX�{�xr��6����Ɵ�,V��Oz�@KK���C3<�������+�G��nbd��pkzD�g���z�ø�RW��β����f�)��$,�b'��<�1;z�?4�~��j�n�%T���b�嵶�ڹ`b}��7�l:5� !i3�5I�>�s9�����)��������({\��q.<x�'������Qqo��g�PW"����O{j��c�5$�T�����y}Cڮ�*栺�� 0���҃#�(Λ3��}�,�r�p�#��<�C5�_Yy#��g�u2s��9�K�񙼄5	�)����]�+N�h�&�ã-akXǉ�TK�K0��(�>�FV�F�LY��w��k�ՠO}]�h삮w�H��'"�!���O�y�P�"��Yfh%�e�5������-?* ���|4�'0]��U�����e2z����]��ൔ�!��]|�a��ʗ׽�Y|�j�<��~f�"���m�W�d�rU?z璛�:�#�K+x�kXG����թu��6k�ׄ��[�۵�u��8ܞ�V�}i4#��^L�^���n��`�����m>�S,�d:��[0�5��N��T�oQ]3jc������X+�qB��vS}F�ZK�a;�C��F�O�1���a�眽�Z���Ys�Y��=,�mUh��p���)�Wї��:���L�\��:M��q���A�Ho���0})֎3B
Q�ּ�4$�>�Z��+��R8��.���;m*\U�ҵ��V�9�a�(�9$�l�X�[y��.u�vẙe��sg�Y�u�K4 �Ӥ�ӄ�U��u�Ƞ���}ba�����+-�X�H=�A�\/F\5�?,�7)jg���7b�M��_�]^0:r��95@��z�� �ćF�l��*����w��Fz��{�^O:O��,U聠�v��R�M�YDE�q��J����[~3�|LD��K�Ҏ �~%%�Ƶ�M�	�/ڈ��*�eè�H̇I����lk)\
�ـe�
���8�o�~"�v'��ĉQ���6������J�]�4.��xg���
�TԗI"�w�����7���Y$V	'P�mz�j6����ab"�����]C�D�%�5k��M�s��}Lp��X�Y)��3��ש�H�K���cm��ʼ��^d����:�0j�&�?=޲���f�5�*ʮX�T���4_GO����r;���B��"�����qg�u���d�����wΥ�w9���Vb��!i���"���m�p����;�sq�HUE5wp�u������f�I�Ɏ�4�kugb�Lk�"��y)66L��*s���C�0C
��O�����O�3dE����Dd'?�jҰ �R/8\%�&5v BK�2�gd���I�J�I,pξ$\��Wz�[��큰hP�D�T���_Ǯ���We@��)����V$ˊ�r�\�ulNP2����F�L�`�8������S%�(�U���-
�O��5�a���>�<ȵ#B����b��}n��u�9B��Ra؃���oE�:��p���4"K6���^0+��D�Ƙ�I�F�w��+Inhx'����g6���}Ufo*��O�x��UzX�ou��&��D�?��H�L�݊�w�zH�
z�}�X��\s�W�>*�[x�t�*c�浽��K'���o�� ��BX��x-T*�j)�Cщ��<�奚��2Gl-��=������.�U����e�c�� 9�.�D�4�֊۫?��`u/[�7��b�̡w�p��g[6xUҨA�$��+V��#G8��Р���4���+V�a��b�i�aQ�I�ϵ��V�����58��m}�p��j&�����j�oлl@����x;/�8'�'�{5E��ϓ���wQ[S�n��,o����,����uF�+j�����m��'�,�J��ë�ܤ�1�%�7}�*o@}�x��m��}���-)��ktc$����e�3�h��y;�$7(X0��j? *{���Az�t�D�]���5� �>�G�Hվ�Sk2������Uam 0<��O`�ŌV��M�������8G	Qn�ت�g>A�W�¥^z�O��n�߿�G�,&q��آ�� p��#lwl�>�b�Ϛ��R��/j��e@ò��C%�<�V���=�:&@<�1HXf9�$m�ѽ�]UM�uC5��7<�#Ej�d�Ҡ���uۨ�q�y�
�����ބ%]�ݫQ�/4�n�ۏ텢�u.��Fѹ1b��CE�c�;�ƱP�w?;��u��L��u'p<]V;�Ġ�u����~+@�~��6�/Kwo����WݤM�m{,5��ؾ�=�G:4�1���u.P���8=x��+�Mnx�EF���<)o�Ly�k���e���s^^B�@՜Y�����0h!Fo����s��o��2Z��i��K	�ͻF�'Xy��S*�Z��*WY�E�1)����;��*Į�hάrAp#��Do�d���%M$T�J���(����o�I|8�g�̶I�RƗ��R��� �#���bU��ty!���/nՁ�*[  ^���{���r@�� �>rf����z�@x_�y.��}�d�ͮ�{f��'� j�4Cf����f~8�%��ҽX�ӟ:�FH;�~ʪQ���w�k�|W
x�ݱk,`�5�����W`\� ��P��BY0b�V�}#&n���ܳ�N&�`����f9�#d�.�� ^҃��p���#n}�ҫ�n��(�)!W�>�F~��
e���tU�ab?x� �g�]���]%u̱(b���hW�8�ԕ������l�r�p�����Ģ��,k��0j�I�C�R�:�k'��	p�����5fu|���d}G�P(�� ?��ߒBJ�N �d�|$1��uM�ל6�����5XKg���|k�4&��^��0t-w�o&�#a��Jؐ8�@��^��a@X��gU��*����m+lc�DSX�{Z�s��Q�T +d�ⷖ�@?9yٚ�^d�Q3�xm������7���xG��+���|&��X�%�v�VR�#�O�bq8���S�[Ϫ$�v�le\�1R��a���M�flAH��ab�������
1����� 5"~~�2�5)�
U^��V#K���i�d��wȍ'�=���xVG]a���?���I�@E���$�New�  ��@���
�cg�]p��^����������*�cF�/�p��{��;%쒽�^�v���}�[��Q )R!�Ls�~�Dǁ�f�Z�n���4��G�5Sl����~�k��L��m$I�<\<��bSCSج�,��*�`�k";��Y���{#�5�م�}�y�Q81���F�Et�t���(�I���CmՏ�`�x2���g��ӆf�',}L�DV�GX�>�s�:��Jm�F��IK�l8�M}����6�Ji�19�啮�
�IR>���!��q��"���݇Pwg̯�Jk�D��(g�hh�;P��z	PF?�S3f$ԑN~��5jB)�z&�p�t'����Vݥ�W�v�)r<�O�6Q��q�&΀��L�Qk�s�J��v��7#���A:��y����Q��*f�-ĝC[�Q�J�c�j`p�䏥V��<"�8ru@�u��u��b�%͔(�7�PuW�}Y֢���i
��_��ry���kG��H���=K,Q�h�i�P�͍� �֨�~0+���� �A�f'H)w�T�����)��dօ!�sc*~��=�Y�ꕘM��eT��̏���^�MTq-w-��E�)H �%�8Y�T%������\�4�6͸��I�Ru��Egp��.B�}����:�EC+��Κ�{,��^#�n~����RuW��Y܄�q��f���D���P�pg��^Qh���a�uM���̕��<�	�T1A�U����0>��.����8�([Ƿ2'^��F�*�`~��?�5�BO�<��cL�n5�}�0����ܑ�4�I�����gJY�K<�_��4K#R'ify��z�K��������7��8�6$
҄�Ԣfx����/cCv�OQh��P��6����%����D������MbmӠR�t��6�#K�ژZ����*�z	�9� ��\��"�#5�W����Ui���0f&�`�Zm����[-ɧ����d�Z{�;��N4��t@P��@tQ�:uO�}���j��T�P��c''�A�]n�i��`���8���Z�9h��UuX�h��OwV#��@+be��!�V�BO��:]d�"*mɴ_c��0�4T�s���y������F��o#:9QJ�G9ظV�G���H��~���b���h�����|�ԙ���v����4��U/a�`�&��!�cB{Fcy�>|4AX;��f:w
Nߐ�Ÿ�;�����3xP,��y��UH��c��i=H����Ê������t��+�oKr�'�f��Ú%=�!����)C��:�ݹ�ȑOՋl���[hW�~�c;�Ċ���~M�x�v�F�+�cpT���v�����n�sX���n���Sl,�)���P	��>�;�5�̷�j���ݴ�:�YBˌ��VEFa��X����D1���[>��Q��%��R��� ��	TaF�~�>P��n��h�8Kz=[���g�"._Qf5���Ҫ� U�i�[:����l�g�d&������~��:3�&�{n���]�-xҏ��> ��9oa1<���~�I+C�Q0)��M�L.�+q#�9 d�fj��]s�|��5�ry�C} �5^�49�C�;�[eB�#��w�N�R����Ӈ�f�Wh�f�fׁ%�r�B��-����
���F��U	I��p��v_	S%��$�)�mc�tB���9�~&�z�<K�-���CPjO!AG.���Oi;�_1\%��PJ]��]2��v>�HA���$5��8m：�%n��<]��y������I��R����,���D�����~���R+
��� $[�+�E��A���s����ypui%h�N����k���8���j�k;a��6�?�)-q�Rky�F0����O�~��CFb���'s?���-|Y��F�R���Mev��~o���ל�h(G5vT�Yȼ.5z 	v�?�v]ã���4{p����,c��*�c[w�	��/�Y�Q�H�'-�^�`�Z�t�Y�`/��n��y+��n���sN����7
�{�]�\��?�QX+����`	�D��C���I���%ڡWkn
���{qJu�r��6J��DT���t xnb�'Hs*&yD���M���$5���5�J������8>Yd���2�|��3�yչ�������(������3}2���@�	��gߣ�ٞ�56�K��
.���/Q��UK�U���3Q#���K:�!/�9s�ϱ���#�����RDH�\D��4�fw�m��[��'��~����3�>�Z�!4_>�Z��F+B�h�j캁�ɒ��B��+9���Vpșh #��r�l ����fPݧ�Y��"�cӁe�_-�d��n!�1�U�e�R~O%����Y��ۅ��Bf�7I�B �IGzd�'aAv�ث�
��QXD%I�KD�Kz�_h�[6>���B	?m'��L���_��L����s�sG-��� t��z3-��@nj��R��i��&��wqco| dٲ�g��� �R>��U����5��8��0����5b��3�/}Pn�Q������A.�����/�3�I	p����A�}�]��j�+$����z���,X# �Ƥ�<��</�����$�r����d���Q�fc(�L�(�1��t�pP�0#��%�w�����B�6]K�гsS>\$RK��[^�ε����Ns�k�rNJ���P�?�V���`���@��j�>�xM�E�|�xV����Z0���n�3�e����s7h��b�ߵ�9$��� �0�qz��F���/@��Xtq�]B���,�X�m���bJ:1/u�xy���Ӟ��Q;%6��8|3L�V^���\����NՍ����[�&緀K
�_x�h{҇ �����N-O�.r���j���iem�5npfH3��&���h���`���A�����e=��K�z����Ǎ>�)��Ǝ������a�W��zL
t���o�`��ь����8	�!W05������ɥ'����N��wIk�%��(K�����2	 /�&��z�YXC��R�U5�m����|06ꎅV7��0irّ��Y/kŷ��֖�Tc�@�Xͫ��� 
̍K�n����$�!���z��~�-c5@���ʂ2�l�Ƨ7��l��)� ��o�e����&_�uC+�Y��O2�'8aȄ�t�HkU��>{���g0�24ߠ*�Aꔶ��gH�f�g��u�wR(���:ɕn�!VP�]��N��d�7Rݡ�{�Ī��oU0�����[l{��|ZmV���/�d:�jZ��vhK�D�=�V����E�\1�]��n4����ːC�9~��>�d�1{n)�0 ��A����[&sR�+*��ZŐ�4D.l�{�Pm�h����<2N�>�\a0#{�H��H�٧/�y2�ݢ�@����[eq�W�S�܍��tR�T��ʓ	=�oe�������}-w�iI8�����6���4w��3vvp��h�������Lig���-�}�@�R�:��rT����X�Nd���ь�NqT}�p%$
������h�� �M�5iQf��Z4�y�*�;#wYj��ٌƐ�����"�g��H�(��m�O�?9�Z3����T��&�=�,�1�·�)sq4��e�Ϝ(#�ĘneC�qeB����������ɵl�`B� `�u�D4 F G=���O� ���C/ٶ6Nd�M5�x^�Ε�|.�s��ǹ[���΂���`��G+��ᰒ�p
�:�^�>d'R�!��}<�<��S$��7�!�\~M�B�
3���!t�X�HM�k+T���z�����0�����8�W@�q|.�A����У��1�_b��� N�|�#-�6?*.d{j�`n����E�I`:��M�R��5K���}@O,ى�H4e�ā��!��Fz����:�������]ý�ȷ�L:��3�|�M�Pfb����l��m��-��B�#@X����RSP8�c{�_3p%�����>H�V��k���k��%���S�ָ�'�*a����%�Q*_Y?}O��|���G*Q҅>֗��+��n}b�{~����]	^��(UC�����k��Z�(��턤��_��U��q����%lQ�<q��e�4`�<�I���9��l�<,�w��n�)�
�r���,�U�[��2mV4�w�sbׅ3��@8M��Y�JNҹ>F��֞1���HГ�a�n���ɥ��IK����3�D��%2��A�/����R��W:W�)��X�O�������H�K���t�.�w�ͽ�Ґ��s7]�~�~��\�Fҟ�ڬ\��\����m�sh�����7nt�K:��N��"
���赏�l��0�V�ˤΘ���Űs�^l���9�^��;-ǝ�~�A��ko�j�k�(�n��0�U�CIF���d�G�h-Y4����{L�.c��:����}IX@��<gQ��ܐ�[�$�m]:w`���	2���1�A3$i�+Xް�?�=�k1}J�������-�:�}���]V'�}H�ơ^��Kk�n<�Ә`z\bd��Qae�M�����9����9�3ʋjh�0��]��m�)[����J�y�n�S$l��gc(���L��=�qw�4lj����,�D�1G<�m�����m���L^���x�zrG��5�k�Џ�P��\���c�WP�/���f_�(l:P'nz-	z�>���6����Po�|��p�� F��xIF��硳3��(�B�j5H>��Qw�����G�x�l&���꙾F����mR.��h�I5�Yy��ŀ
x}�^��W��"m�O�!��4��k��(���}}%oKDk	s[���e��m��-"aݔ\>��i���k&��l�̔ݎV�y�ʠOM��M�;vn��楓+q]��'��p����@��ӯ����fC���8�����_E���Ո\R�=5;[&�	��e��?!���ץUg�4�sx���h�1 ����r1��T�Iϙv�lb����EQs���)aXϸ�<� �%�!�U�iB���I��0�
��B�s N��/�@���	��
k.�7?�<��"�Fֻ�X���b�ձq�Iش�^{�6�`�~��w��H�j����Ć4E�Kx"J�!;?�zZȸe�}����)�c�x�3�$�&I��U���c��W'���I�x��bW��}(>�߯`�-��Epk��i�E ��Ѽe*i���f���k:��))^���g��E:Bzx�rD���|Y#�r5��"�#�t�@���)��=DA�7�����p:bh�!�A��Fb\��^�'���櫩��E���En�2?f
�rk��;κ�2PmB,/�Ҕh?C�-��mh�Xh)MA�[�i_�aU4��Y�C�~��o!>��#rBUg�!a$�"�.k[2�̊�<�Yw�����i�O�H�;}���F_片W���W� I���y,�y54�P�9���2#��k;��*��ף�b6�v�O⦾��KF�}&z�� H�y�#��rH
�C],02K�,�w�d�T�Ji��cGER/�h���Z�pt,�z"�ʂC��r�M�[!G��j{N�w=�4y��P�6�$ߘ���;nlo1��[��j�=Jj�E?>{�	� \5��[i��"!TQ�=��F�ɒ��~֬�KyD�N�֎�^��歕q�I�V�1u����%*B;h�ƟŢ"IzY�=��I�j����ʵ�Eܼ5���wke��*K�hw���������:�f�z�s�����!Zo�[�7�/�/����}�,\p�Y,�2>ǫ�-gT��Jc�2�	��YM���{�Jg�b���%���h+�k�-���;�^���� �tF�M�&28�vO �lk`W��"갭�eک��	f����7��_�!#��>5��Z������o�J��:w�a��%$_��=a���=9����Eȓ�򑲩	Pd�h�<���U|-lV�)t������퐸wT���P[�!ܠG�4��Bށ.L�?��J�d9B�o��4mK�Bh����~=X��8'��٪�u�6��)�A�c`�"����ՠ{������V���0��-���UÕ�Wҁ���xO���|�:�49_�[����}�y�3Y��^jU��;��fWɐ*�	4���Z�u������I�7�2�4�o΃
>�[�������ê�7z6��R�H�ۥ�!���m��o��?
@��6�D�iu�����!nh{��+����6�SE�j/�E�5�۩p]�AYG�1�վz\�"�t���:���6��P��h�usH�.H��ک%�{�0��1��6�-�����.h���t\�����QUV�m�W����-�#�me��4(��
1�D��Q�@��f��6KM�����Թ�3"���hy[B_�Gզk f4J(����s��0��c�ؘg��-�*�������lp����Q��&L�O�b ���;RD�R0KN2,\�q\t�������%�cU�I��to��T�B �Qh�>��o��G�^��<
hI�F���)�p<�HgS��rN݉�HQ�b�f���נ�Q3h�6Z��`���+Η�̩;7�6�g��p'
�]�ޒ����#J-ӵ�#�L3��ML��qd� D	���F��5��{�$3K��+�F,�͓q��L��軍*���}�3�"Z��KZ�ΪW���8iK��`1F@��zs �����866;k��i���4tR:�e'�HD�Z��iJ����&�Y�a��e����,i��h��� ͇v���X�E���?أ�l��<����N��gᦼ�F5RQ1��E�P���o�x��	i3�V�,��k )�,a��1k�A�? u}?jhм��E�\;^y���6/,O3:����=8�5lm���NZRPἦ6�>4G��S%
B:v��9�u�� s,�s�A`�O{��O�*0��ꐆ���o��w�Z�5�`�~x� ]$�@Ҁ籇
T��}���K��eW�=���F��}w�16>�rR����K6)�yt�����o�V"�_he��v��$��%�.@�C������ftH=$�3�2UMHN]��>"�%�L��O3±2ZAJQ�g ���m��0\��`j�;ORDֱϷ)k]�h��Xc#��h�~�G�j�J����R��a=�!kq�o<����� �^�d�^2��$��+ϜR�c�N�W�b�[��3��-��/��b�@i�a7���V�l����v�����x�]��y����O��!�����Y���JXENgw�e'�Y��d�
��3/`�y�v��j<�%�`��`0�5G�ʲ�l��W�?�G�hs�	��f�2b�3���I���p&��A4���4�ß���tz��O�x��߈>�U���A���
O�nGY%�'�^ ����A��u��N���C+H�;�u��S��Is�k
 `��ؠ��?�
OTl�{[�q�V]q�I?�6|�LڗЕ����
����㶌$�5���S��p�"�,��z�&��z��
ݤ���J\�kx��а�/������1�I�����P]M�q�����ց�)˶�}�hK��Bq�h�z�H���lZS��kd�C_È��"�[�xy&�q<�NR]�o����W����|n��J�	c����
ҭN�O��=D�}���PS��?�τ������3T0�ѽR1!im�u���
cF(?k�b�H]qF{�su�'��j�B��K��ؚ�Ix�qt�{2�n�(�d������b���*�4_Ɋ�e�S��]��3��/��Xw%��,{HM��L�,1�,qK�yr�C��F��Z����][�k�,��;P�NxVUu�Π��D)���V2�@��P�m�c��<���������H~!�}F�.߾�q�k�)&��Bb9���=����,{ͭ�N���mL���M��c�0�k�xP��X�#l8jT��č��W�vg�8;1�NMG8�Jt��P{4�+^��s� &a�N��iGR�rN*���=��F�6�./���;nO>q�p�p�|��+	zcz_�r�9���4&�����E�/�MjuG4�����/�z��������_�aqtq%�vl>{ɗE��Էx�Xp���e�'/~��^�u�R	����u���t�zI���v[usB;�$�ؿ.��v�`�I3X�M�ܲ*,�֧O,����H�}"Q+�S �8�����z���')�e�������W��
љJ�����q�uU]��i��1�
�7�t�,�!1���A��������;/8^�g��u�l��YRi�1�K���or:���ʖG�O1�[�)V��1�ŀ;�>?/�I�u]�l�I��a{���_����"Yt�?p�I�m����؍�y%����0Հ�eآ��o�f���T�g��L)�����苻3��j�I��Fo,e9��j�x��t�i��T�_�C����S{~�<M�*K(6E���һ#8�j$��6@sXn+$<����8�N�}x�#�c9�6n�Q5\ch2AWB̜sQq���E.y�t�^�q��m�@�ڒ��I�]%�$�
�+��voF�Pyڌ��^�x�'�gy
�q4�k�hE��yxܴ�)�zPFB]��Wh(\�J}���y���� ��1�2���UƨΉ���L������*��<��_jC���:��뎪��y�$W	�^���"��1��
�z2�J���$��I�S\�dW6�_Vc�eAb�L�Z�'��tT����e��ѵb�µ�y� h�<V�G��4YE�~��cc�XnT[��<�h�9��O-��2]���L��@����E�=@������!�pT�qw)�Rӯ�nG�C��+t�|D�����W�&�{�Y�e�U���{'����3�Q�q��\`ܚ���A^ʭ�GL�=Av/�c�#үP�.w8���*�E���7(@�0{�ˆx���&����z���}�vjGA�<@%��Vf�El���X�����Yz,q�8�W�2o ��rg�P�I���51?x�h/|i-g�����J}��c�#�����`����S�H{��=��KM��3ԙd�u��6�HgU�3A���I8B�"/�a���O#u]d�K�V�~�w�J�Z�LkقU��T�	�����?��?��#3��7�"���F��=+k?��[H��z4*��;�ZnoRčUI\���������%yZx�����̸c��A;�"7���[l����[�L��׽u��wގ )�J%�����M�I��8P��YܒȠ�5�&���RZ���Gͻ2z:���
���n�<s�����e����	�q6��v`#t���m���U���}�7U�b�Vi�k�S��*��냶K�L��kN���Rp��p �4 a����Z�E���]Zh�;j?��]?����suFt�s"粼3.�HlqB`D ���@���~w�̬���1w�
��c+*ǂ��I<�@�'@��[G`K~`F��[��c���]D-Fދ<N��w���H�`"�=ak�Q7���^�:�h��	:�4�M"���.�9�7������K�
��i4%=�P[����C�-�c��m�¤�ħ���馺q�}�^?�շk]�۱��ӿ�+%�%����נ=VΡvko�aJ�����3z�GxWZ���_�<=��бξw����]l�M�Z5s��x�PJ��kϲ�x��8>�6Z��A�]����Cd񴋏Ҥ+6�	��\`�%�*8l��cg}NfعP�*��Ê�}��{Ы���V�%��ZY��ɿ��:��\I"\��P:�({���ô���Ŝn�o�ވ7�g��iZ�}/�e�L��~����I}��Q6�����;=i���s�;��u4e��=�Ol2�.���MnǞ�5O��{���<[W�A������=�X��rM��7�Q�yPw�])D�5�X+2�=���Pm�������Ѡ���Ѫ
�RQ����*�.��C�e,����W$n���F�qv�"��-;�fʇ���7�S���gi�Ѳ���s*c���{�f�N�X�L���|d�D��f�5��H�m�{/�5x�y�A܌���V�=6y^�����_����J���7�42>����Wӌ��K�6y�g�k�if�&f��܎�4���?^���N�ǵ�P.���;U*In���
C�A����9 +k\��C�e�,���n:��֯I_1��r��4PmE�y ����KE���6�T�Uo��\VS}�*���־�մ��[�#9�����q#�0�M�B�j�]�(-�AS&4�(Tb~}��Sg8Ĕm��`s�CEa��d�=Ƞ->��t]��w��^'V2���U	1������f]2�q���9jS��]i�������zX�X��0m���ANs|]Y�l��х،T�4�S_V)�%�n:}(ʚy�adV�Ps�|�h���HO@d���b��0��E�SS����V��B�0����[��0��5���.HU���\�es��X7b	�|P�>T��c�x����{������c��]]42"��)j$L8�K,Tp��A<�Q�
��_�:���aT5��c���~ o�_��M��@����Ea!��>��|+��	7̨�n�7�4�C7��2#�S-��t�c^%��K��� :$`��Y������&	�tfE<ø
O�\��;5��}l�W3�k���I��t���+�q��O7�q>�H:
�x�l�9��E��_�^V�.���dkNIѯ}�[��@�J�:�̧ӕ�2VX��*F��+�%[6�E9����I��Mw����XO��n
��������������ذݴ�������놅Gp�+vd�0����@@���X��1UPPH���ujҝ�t޷�]4/{�OWe8��%��{yW�pW0��ȃ⍖��0/��d{��3qO|G�d���>��Ge����/:��A�ټ:�n��Rɢi�S�=�񻚼h+�|ZC��;�� ��8-Tj±n䙟őA)&ڤ�rK�~��ζT�LŃ1��6K�u�h�;}������ՇFX��w^d/����2��Y����ޚ[���36!�Z�� ;�d��$�\S�6%M�� �I|K����������%�0�	��8f�m��R*I������m��P� �����H�U�0����cW`�Zh_Q'��V\�}(���~���ܑWѶe{�?B��}-m�U�Yq�fnz;�p�qnh�1�������yCmT#b�W����U�$&!U@�f*��[�.j�%�+Q�o{�Ӆ�� 0b��s_�K��sy<b޴��C��C�[p���8q�����n��uw`��MS*�>�"�R�_��M1o���9(�&T�A������<�2��I��ȈRd`ڭ��(�b�a?q@]�j��-!:������*@	q���&�d @�H^���j����<��[n�
�4��OӹŹ���-��?Gr"�!��u���O:����<j�є�4��H<�#�}�/;������͉�C���{ (9>�R0��&�$��9*�捘@ Ib�xI��F3�L�)��iy'�#�l�H�JL�?΍W�^F�9
���S�ʑn��T�u����i��K�-8�5��D�q�Id�F��[%�8���Z��By�O�E�̳�F���}����o�#!ˠ5Q��$������6��p&G"fX���t�vM�DmeNĦݓ@]����\�[?/��l;���E,���z�Y\�5^8�+���c�M#�W�pm0U�wTj�H#�HfJY���V!< ���_d�(�.�@��4� ^��� �űp}��-�CMǵ���X'}�i40����A ��XK<!�R��Y���"Döx<��L��&��D�r.h��U��d֨��#'�eޛA��xTE0%� �Z���.D�a�dD�_�hpw�Q��]Vn'w��^���a�+�g���|�N����5ET^��=׌W,��n�r����,��/��
0���%+��zU�
�G�����/����}kVJj%�C���T�ú�'.#�l#H�J�װ�k36�Ac�~J��Lk�<c��o^�v63s��	�ȃ�+�e����S6%���>\�TW�Ew�(ʣ;���
�븢d��>���Q�JW8(M/p�.��^�f���3��;T��9\��Ui�z�/!�ߢ����>�<����	W?�MuY �F���}���#2�Xtp���hL���zN�S����F�U���c��_J@u�o�\�eM���,Iƭ�ܭq�Fm+�[RYp�f��)F4:�E�i��3��0��`?��
����a^u�-]�ه�������R�z5�N,E��+ݗ�����`��.�"�-��<����0�F\������26�J�1���iU��k��OeR�I4�Ƞk�a�!�:��XbN�*Rf����$D:�j�d�Mv�·K�|��h�~0������l���!�z�<FM`"�Tm�&��q�1�]A�����4�z��C[�P�M�쟊y
����|�?s���Q�޴쵭pJv���G�<;^!֝k�V�z���B)]F�Q��P���	��*���x��R������Y�?��t�4��r0�	FSJzLLBWjE�W�#}31Wxs�zq�j����x�ZN���F�GQ�>�Hh���7t0òv�����o��7���������3Vuww�$M� �W�f�1��GN
�L�)��|+��j����Fq�����5뻒�|��]��m:a�I���\z~���h_� ��F!4M�c��%��v�
m4r��`6SXJU�+aM�.J B��ӷ����3I���}]�rS�`���Bz�A���ֺ���Up�͈V�u���t��wʢ���b#�p�v���j��n��n�z�����#� ë�V:ydU��F�����Ƞ�5g�|�����)��{.�h�\�o���1��+}�H�z���nwι0dY���)i=qDh�Gglo�Д/w�?t� 9d,�C��(<�]�3/�04j-lxB�>≾&q�1�l���vw=&�5w�fx*��p���}k�գ�G�^�#��n�3�+�_���,&oT/�"F���<�Q�c���,8۳T�Y�$b:.-��0_W�U&�,ds�����"���'�n�e�2zH��9��jAr��e�D�}ݐ�ng��q9��:1��EiGÕ�x��8k�Ԧ��[H�"+����Gp5J��*ӗ��;�-�S�����X>�{��!�AE�>'��kz-��ELVs	Fك�*�u��42��Vz(*DZ�;Nڀ�,��9~"zlw�e^[����F`0w{�[���s��Ep�#7��O��kX��R����el5����Y�T���F��ifVL�Z� �>���F�ڥc ��'���ր��V�G�ǩl�l�������B����1dI ����xhx�3K�������<z������\�B3C
Kfne>�_�N$��zb���pz�LT�88'F�A�A`j�P��g�����"�|�^��;F�r1l.�@rMT�#�%ė��B�TCh+"#3�Go�����m��������>���g�c�����E�@��p� '�;jJ��mT�a�jP2m��-6_ƧXp�ZcՀ��@Iza�� %��?�DTڮ�6���mo1���J�@rv��b>xIa����As�Ԋ��rj�.b��O�$u���OX$��� �pwï�qhH�˘ҟe���X��Br/�U�z�;W��UV��i������.E�xbD`���/�~JI�DϞ��DXa����f�'�g0���tlǉ�d@�s�b�P����؄��=�6����}n��C���_����;-�����T����p�3r�c,Pcg`	���辧��:h�3-�A�f��{Z�HnGgv��θ����Yr��v9�8�ſjL�sZ�-�S*����wZ;8O�|� lI5ʧ���g7� �pr*��'*`�ҏ�VCį@k�U�_k���$]���gD�\�b`�|]������|�K�<��V��C�jY����s`�2�Ȗ=t��x+� �n.a�7]U�?Ԡ$����U@8K\��U��ڠC�k�M���P��T�>x��S,��,�8�篸��vh<�c�
vz�y�O8� db���JÊ����F>Do*��׷���4p>�U4�tf��U���|����"w�/
z�֜��W�+�h�)?���n:�}~���y�i�H �rҤ��_gW��ڌ���'4�����Q<��UM��`��U���\�ӹ��a��#��/�!�Q�Gn�K�ow�Mʹ���q�ӧ�>������P�6��D���������n|:��{]��t���H���D�g�ܐ���a�[������΁Д����lj��~�ۺd��M��^ EvV����F$���, 4���Vʤ �ߩ.���{o�:Xd���g������A��x�B%Ym��2Z��a���n�b��}Q\��+���ڹ�"RC^��{@�q�IDu,��kJ�;m�_�K���k�^�jH�?m0跖�b�_�a����k��ɕ]3h�¯XQF����MI�Ί�k뒆 >!z�y��{�qd�(<���=OZ�����+�o�3�F3�z�&Xݪ��s|���ѮWL���9�ߢՏQ��v�]V.���C�O�ZX�����"��q|��<B8��蝱�x�ؙ�"���J~�-�QT�,�}�!*�V�&�����u[���T��<X~R#�Ŵ�);\>U�^.n:f�z���G(�D2�q����<3��{��z.V�2� ��c��iX_ u��D�w�C�t1צ+�fx;t����vgŢ3b�L�>ڛ��OK�ʷ�ΰ��5�ӽ-WbM�CR��nk��;;�f�
���������lo����Asf8ƺ7�����\�ɂuV�{���$Ufv]R�!�l������9m�FJ��HQ��U��^����5��1��^��[Ȯmb*p�H�}N��5�[��Qh믷f��ʈ,�)����e+\�;�܎��m�$�)�2X��%�� 𨵁�~e��<~��9�ۇ�;����<T1��=�т�;����[��n ,��v�IB��8F��f�v�Y�L�+L�y��X��!���_���t���~�O��D�r���s��X�l�n���B}�w�Т�4E����8c���K���j��оX�A9 ���g�5aNdd���,�0uc+mW�C��j�Ӎy�g�T�V�j9�]9�!!�v��XdԎI�{���\������ft%g�TK8e�q�ɑ/�T/-����-���-T�PNu~*��2�s�z�6��z�w�8$��Fk&x�	Nyi����\�>��D�u��3s�0X����P4�b�D^�(FPs�����Rz
M䀆�#c�Lt%��/�����G��
I�m�Ѵ�!*ƫ&�z?7 �2M�lt�l���*xXy�Q-�MWg\/.IҴ"0:ʡ���f�c*@Ӄ�;Ug믆l��:��^`��I��GRj_!��#	b�'s���b}�}cD?{��h��" �R��+ЧN��~=5�=�������&(й���H��=���Gσo�+!���z����|�/6d� t�a�X �'o3�"��bXG��f�V�d��7dO�Y��N��(}�!l��_���<t��n���k�7�;y�~B�s�#�H���ĨN4�����i@��PB ��|)oR#)�x>��\wEV#Nt�Ƥ�x|�x��Q}��ž Q����O�l{��<�,Wʻ�ţ�֒�}̼����4���S�k(#O�?F�N�q���zϋ���=���0���d���L�X��������/��X���H��UrV�M�y�E#[�F&�ϟ�i��Bl���2=E�߲��3�!�ϥ���]4n_զ�6TV�	�G!�K�f/�����ؗ(���n�@������"��K�;�K�?4vF���">b��'�Q�a	��Ztf��L��?b�י5d�a�nb�+̜��V<�߈<��;m�&ADj�s���n�A0c�K���h:�lc��ߝ�ְ܍C��&�@B�)�s� =T&)(�/��y��{�0o���k�ҧ� �/���1�S�yϞ��e׃�SI'fXο�`�`$:ZD�:=���0pomPPl�O�,��9�
uR�S�F�����*��pH��ø�θ{�vڴQeO�\$a$��g?p�Re7�&d���@����Q��p��^�r���?U��6�y�oǨ��@�Zc����Wg����m��<���q9����}�R��]7Qa�#����&�iG�v`)�e9b{��kD�������S�p�O�TP[m���Q�E_e�.�~�N�{��z��R��~3EpRv��ķ�7�ʽ��`~yJ=j9Kq,���r+����{����Q,:�u�QE�7�/���0!�2	Wq,� �Q�/����r�"���Ӟ+��V���Q�~�!q�j�B�ɸ��������g_��etm��S��c���2LDȄ����k2�Y�BӼ��{1b�p�8@.�Gȍ�� (�����d���,�4���n��(ġ��J��`�.nA���[G�^g;z�b�������T���;om���d�T�|R�Ԟ̯��k�Q�rCe�V�N�����/;ص*cC�aA/�X�2�P�s�=N[I}u�� �p�뾞p!E��~v�vK	��|n�<�V�+c���J��V1;��R� ��C	�@�z�n-�i��~�]�R�}t ��q������W�y��׎य़X���٠hv5��Hޱa�$�hVi�q�#x���pG�ӱ�\a��fݠc�a�EY;�8��J�i	8^w�d����������l�^�:r�h������ù�� �7bn_)uF���ޖ�����A���6�fv�*?bsR�~H��2�%�^'��[�	Re�v�wjf�g��#�aR桿'gT�A"�u�Ĵ����t-N�w�[^5��5�)H��d�ovQ)��;�
ix����O�#���������u�����a�ޫ�5vF�ԫ	ݼQ���h��}�/ت��@�<d=z0��h��ym��ޓ�Uh]J���a��
1���᪉����C�#_�d�K��]��W�eDkZ)p��'�7.���������p�[�����w�E�^y_���iqժؤ���T�U�3n�Цpjm�m�.��@d�G��i��~�Lc{t�G_=�78Η��;�7�<S��yl��̂V��BNl�c( q8���#߆�\�x����DFG����K�}�jj=ǃ�E��Z�9���^���&XTυoY��hqb�(�:�Y�X�^�Z�Q�dI*� wș(�X��Mԫ�So��-"��Y_Q�$��3$�n_`͏uI��W�3^s!�i�8�}��8�VΧzݹ��XJ���+D6��5a���sWwi_ږ <��f��B�KLbk�T$)?����[�ǚa@U����(��=��|�Z=���@�>YpE<��",7׶�nKa�J��YR;��O���ލht�3�M��x+5��)���^jcs}�{�Ð��,X�'���FO,�RkT�@B�*��5\�';�eu�99j/��8��Pt>�DV�����/��`n���i��*�vfц����,t���qUK��U���\*�@����1p}�C���f&e�)խ��DuJ�x�t�6fr!��n�Z�p�`&X*_�.��5�rX�D���.2��+ ��9�č�jaM�4y�i], ���2�1���;�<U��$N\��\Y��Y�ʠ��.��v��>�O��x@�?_�O0�M��8��"!��{D�p�Ư0�R7�}�-�J�:����A��!r�.6�ڒ|��8�Q��6;�_��c�9cC�����0��-�^U�	]��CE�����M���K�C�R�����m����y�M�w�T�����Ra��T�gŽG�cl �E^�CL۔9�В���ܾ��x�jV�AS��#�C��m���T����d�z�7h��:��Xo[�Vݲ+G�	��2V����F��e���&X{����o��}����
�e����^���o� �	��5�4�}�V	�{e|�D�$j��9�|&�!�t�~���l��B�C�9��e��"@+ɖ��.�-
$�&X���,��^���q.�:/;�9��Cܻ���u]��*��r�>�`P�:�ʎ &S#C=�E��;v��1�o��V�(��V���z(C���F�4U���ㅵ��z����et�x�S�2c�;P�ė�*-�_b�_Y�m�kN��*虩fR��i��𝕳�����@M�ĘS]�i�j�r�n���Y�,�d>��0�an����i��4��Q����^v_ no�!�!���eL�-�mgۗ�+%�:�]�[��.�ɦ�GЌg�U��h�C�[\���v����!>RO5�6�.`�M!�%����i����ƨZ4:u�0W����Eo:��n�` ˰f8k׆�?g]L.9�T���;��G�o��+���fýv]�EY�]�<��З軻�~�}�!���=o��ƅ��X����`du\���<����*r��Ƌ�u�~�zv��s�x��� �2���+E��<�B�K!;�W�| 0�z=Df��G��Y���Dj�2����{`C��bރ�>�g�����WKsi�H��q<_���+B7Î��hr6�1=�e3�y�ս�������q,��K�(�_��ֲ��D#$3~ofɒ���2���l���1Oo��6R�,���=�0� 1���&c-;J���<�5c�D�z��1u{���m3Q�(H
 �m:/�Q�]���B��>g���K��:��µX�� yL�S��IC����
æ���䤽�X� g�Sί�ui-.���9j�܆P������ӑ0���(�����@n��}�l}>�	�~a��Gxg�=�d��o(wT��pl�#I���b��$��2�����$�a���^��!~8�5a����X;�Vw�V��"��� .������6�u)�^���8%"ą����|�/��~�g�%�����zh���#��]�}ZN7�C��,Fz��ʢZ��V��o��<~�'�#`�O��߻*��f}�"=�~k�Ơ��]�啻�}8z�����6i�!�Wjm�H8
��q~�@]?�����I�4l�}��Ȓ��~>p�F&!j��`��Ijg1Î�2
��6�3�.��k���B(bU�-_q�K�.BO�*N)˧op�����@�Y?ޗl�6�9��<m�Z��F��!���qk�)Os�8m]�i��J�KN+w��!�}���& 3	"�bF�"U�*9J]���;�\��&�g�퍥�M�Q��®q�]��y���9���|�~�o�Rj��|�����8�;2��:�eDo6���)�e�[iC���$�(�ҫEs)FA�J]��=������A4P'���N��B�_c��*@�����j���iHb���]���؆�ihOf��R�zt� q��t�O#���x�bkG!^���~��gK:d�
�q������N��1邆�`�i�Rl�骖����)X����6��n��H(�T81�%�/N�N���V�ȧ!���dD�dL����b�j3c�#�Z�)�&8�Y�tմòP��6�hJ�W'29�41ɣm3ٞ����:�7�\2��w��:��û�7K#FQ
B��nb�d/���aL��/ H�?��(���y=O����/�'{�0+��[�ϼK��j�֌e�m�Q�@:?��f�S����A�Fuk�$�ur/����ĸ�(��ugzyWdh+��g~&�6T�r2��%=Z)/�����}W�hIM����	�Xm���'�O�=�.�nڌ  OP����&Ũ��UY7!���'"�P�D����0va|^�1{�ʒ��\��m���r-˩�	�H6v� *	g3�j:�P&͓���3ǒ�p�ѥ��?���Ds�F��*��vgf�,�ZQ0i��r­�eW��ܻd b7x���$���dj.��I:[����O��a؝^�l��w���b+#�Rr���W��`�����Q�"�ce7G��E5 OD���P?9��A��~.O�:��\�V����(�x&�Qf@���Rn�`x��ҋ���u�̱��E�Cr+4B��u�����&-�m�1�b�f�ób�=�0�S&x��K����P�>�F���Tj��X-<��GP�P�A6�!�1�x�̸ye �k���Esw��e��-_��H�\��Q�T�����H��^��#(R�q)zQGl+O���U�X���$8d���F�Z�����-/�X^k�nձ�����΍��j�����ʦ$k�f���9	���jeMJ�-#B�'I�O��3� Vb�}M����|�y&s���́uy�2�
ܩ���'՝j��b�4�sE��[���
��yo�-��U*5+����t%(�b���lY`�������K�1�)G����AJ��/0��Z�b�����3� }VV����4 ��Ŀ�(���ɤ���x����My^W>ԮPN�ɉߋ�í�# ��@���*�Gl��bQ@�[ntg����O�D��V*��0=q��N�ڕ�����^ޱƦ��(\�֐jnȺ�(���8�f˿����_�X[m)x%Gi���B9f�2Hƕ�L��d�'@��~�?��Ɠz^�{���(��u�S�şp��P��ɝi�����N1�H�D�:�U�b���VL�qy}k�&7���e|��QZ�mkD����p�[��~���!��/U��ܮ��PUg&���moi��t���(���}?;���u����Ei�-D����'s�f���/����ζ������;�I��6?&1M��(3���q��Y;��e�lh߫�g\!�p�)(e�N<��������:˼�)�,p$�VȂ�*�I��H@Y�A"��nX���i�3?/�:����P�<����'��z�?��;#O��K'V���tjv9N���8C\v��i���r��+.dĒz�-ȕrωSF�9�SG�hA���ؙ��x4��z�|Z���\7R��p̍�=���d��Ҧ%86k��fv�f�ݬc":B���Ƅ4\<m��0��]wTI�hG�l}D�t��Y�P*����^�m���Фc��bӧP跌aCҝ������לճ2�����Ҽ��)���U�kWkwC�`	�_�RH�jw��͝pX�dp28�51��aʰF�ߞ��(��wu�j��`!�	���AhJ��_���o��-����#%��<sg��LfoIG�Yv�zH�����C��Z^]�^���V��׮^+.����ꭷ4��usD2��g_���w�=�-+{���'���F��Z'Czt����t��n�����I-�H4�_��**>�ԧ��j|B�3�xȌ�7�u�`��F&<){J�Qg���y�C1Y�G�aHI�\7ϓI�
eV��<�-*S���?�{߮��ɳ��S���q	���Q[�r-~֕a��M�H"�ǭ�Z��zk�mԀ���H���q�&���)�1���|u���[q_���e��j��sՁ�XΥ���t�_��߶۬Ti�ߟL�e�h딊WiD/{� �w�ض� �̱|P�m� 'rt�o#	���Z�	m�BTЖ�	5'���T٩�;Pv�����ت�건�2���� ������ŞL��%R�"�i<�pNA���]bv�%�,+�r"'x�ߙ��ۡ�����y��/�����|J�.wT�'�G	ٜ�����5��3V��z&#_�a��,�W��$+��x*dw���J����=XZ+ƅP%-<om�Gc��_u��t���P�&ы�iܦ�3"O`���59�&�ϭ81�n�H����T���
8���5V�!�/;]�jF�w^Gel^#�đ�R
i����S���axN����	���]�X���Q⯉��u�4u>ba�O��s`�J�}�g�Ӕiާ%�9gD��fc���|���7ӄukk��R�l�V�|=}u���w�t�;�����dY@4�`��d;al֮��i�i$]����:�s�'���k��z�T���-�W���K珵֗pbi�5�����;������LJ��m|m�m�zG�� aѪ%���hܾ��칩Y��g;�������_��e��-`;�2~�g���d\�W�̬+?61����r�t���M~c�F�8vr�q�_��v���:��{k����\.:�������v�%�?�x��\���V.��[���s��s�z�c+7E�eM@e�i�����ԗ�.�ݖ�20"�~��p<S�0;-�Dr�᫪/�+$�@�
�ExjX��͇4����Lэ~ݜ-���}i^@X%L�9����q��� =�D������o�T��M_A}Ν�h�>*jqͶ�Ni]ߺ���z����9�"�1>|^�׬�S���,���4n��c_��i�l�ˏ!5Nm��WU^��R��>�e�`꽑r�4Gmj�`+���*����03��Lȼe�c�B�h1,���F�qF�y��=a\d3r?����}��?�8�cQ ��P���Y(/�kI= �C�d�eTsב��}	\�}>��#�e���!xM�&:O]=�<m�wJ|��h��@���D�:��.�*������<��p�T�������u�& �c!�;�����P�FF3���}���j�
4u��q�)�`r��}����~!��hU�ve�i�r�>Gh�����(j�;N���n�s�N/b v�;a3��H��v��0N�:�̛��"����Ld2?ߧN�a*眩�A�� �mnUu�)���"┭�:#p�� �퉿<���*�uZ/���,��<��vΒ�6��8�Wy����k1�f'����f 0{�x
�Q�b,����)/"2��ӆ�}ps,��CtJC3ڥ�[�q�R�� L��<�C�U�3;�43�DD��~���|o��g�d������Bܸ�N�a����;�� �?�Jl���X����a��|�"$�ͦ-`¼�-�{�����b�C5�0˸�ς>sٖ����4�P���[*�ߍ����o�'�Ȫ�cH��V��Td�V&Li�� ��zCS�To��¿�i,R#t�K'����(���N���9��xZ��2�N��/�9�viu����
8�����(l;L��G@���n5���q�3_]WW�)���ka]���Oo+�:�����M}L�>�$�Vu4+*!~�{/t�Mq^4�]��r?a�ߘy��'�t�|
^%'*U ���غX�d���+�07�N@Rѡ�=K�N?�>&�t��<��,��hۗ{�\���I������@��r'� �io*tp���Ie�>��@�5ͥq��V`�&ǩ.�T��VR@�]�)��	x�B9nX�j�;������r��� �%�E��E��e���0%����LC�gA�&�[f�g:��E����ܘ� x?�,=��� �&�}����k[�h3�"8�G���wg�Ѷ�S�5N]��UGP*\���[�2���*���P�?S]^��G^y3U�a����T�UG�n�qёW���|D7DܞNz�X��ӱ�a5oK߫�9�������UdN���;j$n�>4���Z� cZ�}_Q��[�l���0<��#�c��-A{�bX��ď'�服 T���������o�H�xJl�kd� ��_[��*@Z�@3����&I2pL}lG'�/�,�l4�K[���=Z��O8��j��/G}��F������#_�����Mo� �J�H�B�!@�n��{�ڲH���i�����!����?����]i{6H�f����<k�1c1�W{��E$=D����d��?�{�f���J_�>$��oqh?�3BM[��&	��mj�֞�p�{S�#d�s���E�c/m�[
e�cܑc_ˍwq,�h��ZrĞa���ߠNp:
uj�Yb��*��y�yC��|Ѭ�`+�#�gy{��[.Kr︿R��q��t&��(ȞU�b+���r�n?�k�c�¯��9'����˶�b���0hs]�>��K�mXHo�;|�SIꄱC矜쁁���.�~��G�	��_�f���0�e��Cd�k_|�+�c�? |c�}�6Y���~o�lFe'��
�"����`�0�}|�hv�A$��-|alZoM������뾬�B�����ݷU|C���P���g*����#i��C��뎰ح)�qLs�Şj_{�(0MS����
������˔�U$�l!|�-�]��cY�X/ɒ[�CWJK�f�� �~�ˀu������>M͎��N��or.I`�LePtd5�F����/�q8�Tj���?T�n��
��B�-k�( `����25�̍U����^�L�,�9���_U���'��[��3�o˼�nC��C�K~M��R���E�a��f/�>>���+���f��؜��:�F��[\�k5�������?NU�&�)q�W�[,�R��\G��*k��1�q�@�l�>�H0H��;�ƻI&�WUN6bRU�����:�6A�P��U���#���p�1yȇ��A'�aO(qN����`�0y������I'6��3{*�؅K	HékhF]2�,�g��=T���n=Il�@�`�0��D^�s��Կ��o%p{i9;���!U�[��T�PGb	�4�|�&D?��К��I5D�]�L;�de3������D��3�z�6b?��/z�f�ǉ�UHQ���1�U0�T�����N��r������;����`�8m��,E8Xg M���,4�7��[}n�R.�:�������)����:��)��l��z̈́��<+#N
]��7z큋
��B8�(d_�6���lǃBC��W�Q��s�����PsMG���^�0�<�	-!�/�YV~d�S�o�6�r��\��5:#7����SMC�:���#F����}��%i��w'�fTlY��͇���
_>���H����sDh�Ƈd�o�_G1��IȬ�W�ń�\����G.i���ot�?Mcre����ZC];u�n~��f�ҿ����|=��H�Ų�۸ҢhK�����0۲�#2�4\�l�v,]K$V[��S��t-X�2� ��qj�%�V���c�D�ڈ���z8ƛ�ޫw*��_�0���n�CQ��%�3w��cz.��0���j2'd��s����~U�0��v������N���n)�Q��gEG�N��E�
?�\0�D������ 4B��;��_�
M?<�`
T��t�S�|�n�'D�����t N�Fk�b��7(G�|���1%��<�3�.������bVZ�X_c�����RB�
�������F�*����M�^^fk�`t�ep��%`�&XV=B���>�.<i,롷�l�k?g��'(E��5w"m� �}���S��l��!�K	�a��y�<�ҩ".��{]��=3 S?���Mńļ����መ�#�*�����K����w?N���zK�3F'���/#iє�hi���E"�v��l:m-��8�?���Q�@3o���b,7P�o��O��?����:�����Ǝ�Z� ��BWt�d�,��"Of�R�V�q�ˢt�l�yL�$C&�G����
��XM���+�����%�=A�2ܾ�At֫��������@���᥹HgA�	'["�6�e�5�̵g���87��w��F1o�L*�D�M�c#��|C׿XE6�q���;��@C��qK�q׍�`@%�rFJv��lk���`;�u�V�H2��П27�W�Ҫ��JF隵�l3��&|B���@T��i����|(W����(�݊��|!�84��S����[~3w��Pɚy�V^xث�k?�>��2*��a,pΔ�����^Qn-q�d�,bMܘPx)�gP�wt����r=���]1�!& � �k���	r�}عѿ��C�x�87l�{&���n�	ީ��������c7-e��,%�w�|4�:[����ۧoK�I�V(~b8S��r��x�L5JxV�2�������N��lYטW�u�������E�U�ߖ�Ƹ!	x���*^Ĩ��������1� T�?J�l�4Ou�m%>����*������Ֆ�hG�}	�:O`�!Q���*|�vl��B��}V6Xa)삌�`����u���T�\��)�Q����m��қ #����s@HR�ϋM>i��y���yĖ6T/�;2����JJ͎�y'�)�(@} ��Pۆb�$��ȼ�ՠ���A�����	s�[~�g�ѫH5�/tK.����b�B3���)��Gv��(������I��%��5 z{�Jm��9��B����" !�;FK �؀��p�C�ݮ��-����O.^���9i_@^<n��ޮ��w��I�MvV����6���:�[$D�"��=B�r�F)�}�-���҈n)t�p��\ei<�׃�͉���;��&!�}�n�V.��zz(@�V����@C<?s��~��{��v[�\E�b�e�n��c\�c��u@4�M���� ;F
"��<���q!����`��p�t���p�`#�,U}j0[��л)Ga+늼_[G�GH�
Bm�������ԟ���9\y%��V�Ջ�#��5�����\6U�Q��w�T}B�迧�_t��ia�Ml.��/�-:C�/��5����G0��X]n�&�i�fqxpqK�8�_�n��H���n��|�+���~i~�l/���V4K�g��I���~��o�F�O7MU��������z����%n1�LYw�^U��0��4��J��?�b�1��hgA�%@e�&��(T��?�~�-܏k�����l�Tѓ�?��k�~�&|��	$���s��R�G]�S�.E�%�_v*sl1T�$o�'�C�܍X<r۠����xC�z�«�v�.l�N�>�o����=��28�&� ̷�?6Zt��F���6n>��b�Fa��h�����R�?(3L	�s�:���L��ԊEqa2[ʍ�ci���7�&���'�o	�.�.1N�Mi���2�/!a�*��?�u�?�@�<��,��3��u���'>�*Qo�y_뢵�!Y�Ĵ���{v�̉Ѧ�fzb���[�n�fғ�L�~-I��$$~�#���R�lu�)*sl٩�rЩ���d�D�1�eμe 	Sz��,櫐e�>�1�]�͉];N�=��/�4����\��ͯ_�uJ}p�^%�T�����:>Fm����t=�;lS8~UTcH��[U�TTn��(�m��kt�r��3
�! ^^Ԁ�lP�A�;2��r�v���T�R�*�E� 	�,3��To��1�I��ѓ{�%_�2��bL@M�BM	u7p	!�GL���hmDiH]��,Ņ�A%Yv��\m_۬�#��pk����}U`H�	I�&��8���z x����.��=�}*,=�����2�Ѯ��?���|���2���(��B��Ƣ�zZ�����keƇS�����m\���h6G�W�؄��˂_
GQ�&�m���Bϓ�{O���
?�TM �6�X��@�� ��Q�vy�� "QO�4=z�I��^W/p�8sY�L̢k�FCT�g/��O%3��)]�xw��y��c�K�"�ZE�#��y(!o�k5Ex�O��_q�^�3{�����0�>+Y}��P4b,��u!�����0f]�>q)�ӫ;pī)�G᳞�����y���q �����yݕ��� xAp�y�//��q���L��tDYd�F/��$�8�{�`�߃��/������ˬg��	#���#��s 8�,��k�W�ޝ\���u�ܚmݔx�i�u�?2C�ruUی�oK-Smp�q�p��d�L+S��,~$�n�1ο�pT���!}�Ж�ƶS��㎳�}�k�o��[F��,�m��V�)N$��FsR��??x�FG=if�c�#+`�����E[n'���{�����y�Ϗ��SִL�����#�:�E�o^�WA��Z�c{�Z�:������՟�,����!oe�����mt�Ҭ��/�l��id���E-��|e���:Y����-�[~}+q��G��r�Pc��:�h�t)��Q�0�r����4?.K`er�����] �jl�C������\�MՇ��&�Ss.z��=�qH �F_�ܨR�x|�~��c��#�A�W��%�����ՙ%r���4��%\S��zR+�j���&�*�*�zaG�I�rx	U ���T��o�z�gr�����`+2 nv�k��seH8nxW0S7���#�3���O�����
x�Q��z��.���bL���:3������2[�:�aH+�B���2�H��>�[
���6�۟���Y���7\�_��w)N�b4��i���_�}�}��bV�D�f��	3�EZ��&�8*O��n� �!�)���H�w�>���t����S�
A�:
�N���S�~RO�56�P]��7+Ep;��T@�����$|�
V��ʬ��d$
b�q� ��m`7�;�6?фR���.�� �t�Ԕ�W�ɩx�eLTU	���PU�ݦ�ѼC�]�s^�����bK)�o�I�I�+x��ES0�2����θ:�/���D�]�4uH�6��u��R������r�y���vi�>��d�y�O7���A��s��6R�����R��J�I���~q�F4+�Bgk���Ja2���#C}�� +R��dO�:`���,s�Á�R�m���}��0��w}�+�W!O/u�Z�/��1�V��򘂕����VB-��x,���p���0�[T�}\�*Xؠ�=%(j��6�	�	'��K�����������a�-�>Ө��0��^E�ip=v�1L�ά��u�ս]�}V_����Wt�:+f.�,�K�LL�`z�tdG�[��4����^w�����+�kO�A�Ј�`I��	KNG1���YO>gZ`TR�}�})�m07��|}'6�2��Pp���gk�V-O��Q���YW���`+(#��ݎ�C�wھȑp�s]wJ,:��}zV�`ŷ߻j�j��V��E��N���\�*b��[16�%����.5H��n����J?ѱ+E�˻�O/�!F�(!�	f7�A��U�?�w4�� /�s�Z��ˤ�3P1#v�� ��+�E�E�bA<�=�#@��ٻ��^���ϸ��q�s2�^gJ��8 �����E
�[��,P��ۦ�;~��}uN-���UV�dRW�l;r@�~ 8����O͆i(�U|�e���3�4py��97��_H+h&TU
�+�ϵ<�{N��U�0<�QB����	��6,�J�<��vu����e�����.�T�b�1z=d��X�n:�B��>��݊P<�u"V�������O��Ra!Ƹ"���otK���~�R��d����fAѸTQ,eY��3}Ws�Թ�*��C���&��2�(T--�v���ɝpD/�$������'|BT��{d3�e�n�Y�x�'�;��|�r]����{�;�%�@�=@!���.�|���xoI+��wb��o��
O��s)��M��K{8���^ӣ�-A�����X`��*ث�x��ی{����=����/�f�R%b!Y������L�H������wv�de��^� l��/��Y���l���g&W��a����+���Eb�Ծ�J�	9Zb�Ȓ�K��?���20�7��F'���Qj(����k���<��=�|03J5eשj6� ͹�]���H*W=�,1�4��s2�j����Z�n�Z~�8T�u�����|�Q�C����T	9��\ƥ���r)�/p�RiVإ�i�3@��Œ���E0�����ݐ�RmQ@d���ق&�A#c��5��%'�-e��\�hz�;ڝ^�h��3G��n���`��0����U����>0��$U��9�^�͈��均�r���|���*�����\g��z&�����{���$�Y��M���f�.'d���[�2jF�I�m�B�TS�'�b�z*�Bhx9<\�	���2���:��!2�ܶ��b��"�C1q�Q�� ʜ�a3�߯W<�r��R�X� �kт��Cz.F��M���*G�A����i�]���&O$� �v.5�R_d��,�5���r��L�F��5�����=� $:W����4UUBX��ɽ
��I�.w��@�h^X�<���S�+�]�>!�Gn�
!����)����HV\R5uF���3R%!�x5O��W}k�M��4Y*��,f�����13��\��)����We�l0FAQ��CX�mB��7NO5 <�T� � )����`Ɓn�ƍq��{_g4)75�}b#:���:y�����N�z0؟��኏It��0�A�x��4�H�#��{=4�Y!��	]��۔�����#�K���3�zm�y*vHb�@̝0���&G,�F�ܰ�����8tq��e�����}2�*��Po�4���9�t��v��sJ�ل6��d7Mcb�v�LQ����F^�p��充��?�GG����A���O�ǳN����g�V�Y�V����k\�h�!��c����dD�)�����h&�Ǭ@��f�y���ͮ�VSv$
�*��/�z돉/=\�RhZ�v���%��D����8��%���'q�^]�Y��̱�z�ǽpO�zs�3Uzs�.��9vR��Ug'�����"��J���:*xK�G���1ͭ��u��/�_��^Ǿ(�>2�!�H� /jOt"{�����>���z���������^\)�ƨ�!(=�c+V�g�@ً�����r�I톗bS���n�9��]�?K�J֦'=C~�������{�ӱ�>�V�:JƉ>vI�9hĄ����su��B쀍`��V,?ö�pG�K���%]�&z��U�.�b��i8:�ho�wS�l6[E�Ж���-�c�����<�m{_W��Z����]~p�:H3|�b͏���v��6SƤ�����P^��?�c0�-av^'Rd��!��`P��<	ʼoTC�T>M�X8�5=����^[���8�v���|���M��s�������s�'��^��>�񏺹�s�;�,� W��B��^�D;����X�Ի�_�"��������\?@D
��pBU�Z��j��K��l�& ;RE%��):�����������z�A����k;��g>�����c3�&�z�p~ߒ7�ТqaoUڙ�RAi�j�|(�`����	,PU������p�=_��� F���ju3�b�����#$�m��=?��(�z�{Ե����k�'9E�mmx�R��(��|
�1Oҧ����Ѕ��]����P��� �P!Vӿ+!c�IXj�}vG����b��#å��<�8l�m�i0Xb�K�%��B�Q���O2"s�����ڢ�X�Dx;^����i�&�m�([q{� � �ڲ�G�!���˗�+'Z$�}q�1���@0_����X�UO٧ӓjs�E?M�T+4W�1{��*2U8�H���[j�QC�gpQ�=���h��̫<r�#���	KU���W|�J�D�$���E����M�~j�@	~��=Q�P# ���*��x`Y�����yχ�UO�9���b�j�|��/X	�j?0��.��`Q1�?�_I�Je�{�`-�� �Y�s����B�D͞�f%��bli��9�	�Ke!��[6�|�v��ms>uDߑNcI_I%MF�/~`==m��T�BJ	���H�������s�?�y��F� ���0�;�3��@�X�JJ ���F�VQ'�3}���
�/��e5u�V���g����a��U�F��-ȉbs��uyށ�R��/�/`ځ��~��$i��� ��� ��LE"`��)�e0^u8,����(�<	��(�%'��?aG��ңȭ�j�����Z�9<�5�pυM�ŉ����SH]��G��)d;����d�|H�ФAI43�%�O���q��i��NL(4��B�IP���$�sD�Q(ow�L 7��D��OF8	�
9��r|��y��j�����*�ி������ B1Ċñ��'���i��"�x��[�A�ꏹn�X��4�(,��bcS���y�:���ſ��-�p��u��M $�re챖]f�)�x�|e��fIZ�UC`��o�n���Ȥ6�*���i0^����%�ύ.���zſ-۸5o3����%��1�'�&[��K}!͐����:X��pzW�2 �,��?�-{-����l됩�v���D�g��i�t9� �D
�Ɓ�#�%a�D��*Ƨ;c^q�E��i߼L��$��z���YC�FJ2$V���f<����k��+��d�|�m��Ԑ'��^m���J)uą9p�r�Ԁ���	)zщ����Z�"uYT�BI@��TiIlĘ/"ֆ��P��(+3��$�����A�q�#�Q*Z춽�9VP��r�~*cf�Δ�m���Ľ9͈�=�����+}ǘ	s��"xg���������=pmk}b��pcw|(�iQG{�0��r��!�{t��cZ#%����a�`���FA�,��`���N�pt�����g��=�G#�_�o�����}`�6b�g��7�c٫�N��G����ѳܨ��w�4^�/f�����Q>N f����^�ED�;���ibvK�Z׻�oO���O/%�]9��.I�=��g�^���͌�t�1�t`-�����a��=��q�v=I/jՉ����B0�����=ZW��D|u1r��9	���*�J�t�\�hˋ�T,�&��/W ���r"��yԘ7H�L�I]E w��J7Y��3I��.~�R[�\�^V�:����v�,�ݭ����ueD����ap|�,��c9e\*+��?�<�ƒ�����髐�&�2�A(�����}b��VDȣ�׶���M!�����+ Rϣy ȓ] YuR"x�q�R[�9���:*'#<B�_� ���	r
9�d��O�ڞ�R`���(�z�R�ގ�^���I��)QW�K��f�� s�T�q�Q�t���ta�Sz��3���b�`��Z��Ƽ�X��T�5��S�����f")@5M�bl���C�Q@6�0 g�@����zXT��*uG�W�Y���'�Q�l�W��.�y��	�|<ؿӔ�3��;L�Eq�[
�'��p����5�Hf�NV��Ck��L�}����YQ�˹�0KёXs.��?���H��'�� Ј^�>`��͸(��Sِ��Z�m\����9�\1��&%n�R�m��-�-��0a�f6�� FR>�4��t��R��˃�Z���9w� D�
����<ey���%�(+YT�z�Ս��	{����ԫ�!�7�e�軫��g#�����K��x��xy�p�Z|��9�8e�8��26?Nn���jh8��L�����gң��`�o���sh�[�U�^c,�싷�N�+�Fp�Y:�#���Y��Ң���[B�@ʯ�|a,>��J�]zݽ&U?ќ�_�_&baw$��*�x~-7X�8j�^e��#���E��!��ң�ga�o�:����_-�V�`&m��)]��S�UO�R텓B�`�P�34�E�+�A|�Ƭ̢��Y�Қ��p��#�H�T��d�L���X���
#�]��^[+35�%
�}YD{e}5�!�D�����9�!� �]�>��C--r�UL�z�|�p3[e��r�2��P"/�π��j��x�e\�%�ϐ��F�k����'S�`�il�:r^�[��,���I�{���1�)���s&��CiW����x�����'R�P�M���D���Y
�"IK"��7��5ե�DxM�S�������R<�d#�K����u���r�:xɏ�����weW����@�2tY���[�	i��<����?��s q �0�@Ƶ���JZ��qUIV�ta,hgi)��ȃ�+I�p�hSHtO۴�E`�����q�pʪ���)T0�����~{~�\K�y�!�w6���@
S�� �.�	�ü��hV�s&Ń����O��­�*� $L%��>��v���f<`�Ċ�ƧS�m�g��/�Spb��gj|"�)r�m����<o��qK�!G�E��و�@�p����@3M �J��I� ��D!/n7����ּ�����p؛[�������~��琌�9P�j��&�(�_��9EvV�I�=�y�o�a����F웦�t��<׭Ŵ�jz�@j�,�r�ʀ�}�?��%t��@�ƫ��_��g�Y�T����Tt��Kĳ��&�P,["��
�&A�M����,���� �x�:�{����;SD���<��E������P�� n���FiNz�)Im�&\>��@���� S�����H괈J�b'����<ɖ�ڽړW8D� ��(}�dʉK	)�؎9}�M/�[y� �Gd��P"!�w	�2�������@7gt1����xD���'�Ax���;� ����c.�x�$-rk�~'�XKq����"�5
��/��T�¨)皥I����Wy���B�B{I@')[�7oj�RƇ��~�;��2s�l�h<�㿽g����mg%�M�Է<�h����ߥf#�U����Uà��x!�}=!���xP�6��#�hށֶ�z+����ԋ�e��x@	X�*Z�(��^�1�@3b"\;�!cХG�FSQB���ũ�J��w�1�4�=ja ���d�¹lab����q C2O�/��AC��V�_*�
W[�T5��ۯa�[����=L�ͩRY��`-����W5'���|������/�"�������S�y�"�Y���w�py�^q��~z�S+��t&$���Lp5wo*�~��l�&�#�of�0��>3H�^
5b����p�ڸ;O�!�!��!R��48�8ÆxK��H��iӛ�!��Ƀ
�!������m��:*�W`�?ԙC"��?#Ka$��ӳv�$֞��X�y���ӄ�ɟ��̉. ��0�×�<\cb�
�eO��Ù���Sd?0�澕\K�@1�fMT-\��9��n�MW�.�P+G�a�9�7���p?MQ!���!�-�qp)&�Cz	�O\�����T�d=���ej͞�9	"G����>ʼ�	�!���^��^��0c�|}����黈��Hf�Xȣ�΍̤�3Vҡq������P�������bg/�O�?�p˄\���Y�m��`9�*�tӌC?b2Y�Gwy����m��[^�(��	�8��*>*Э�r�؞T�jE��$
x�B��w��t0Ԙ
Ĵsk�t���5�;O~�j|������
�������b�BӻH�`��#f�O��=�u6��Ғz���b��C| ao��
����bB۟����Ev�v��y>1�K�e�Q�Z����������׍^T^�=��i�vG�!7��/�i���o ��$���0@�M��b f@�򋝺d���~瘀�#�ǝ,����s æ�X�(�EQ����´]�:�Ǣ�X�[�Aӹ�32
��1�d� ,��� 	DՈ.�d��@����B{C �)�o+`���%}F�Ĭ��,KLM�mdV�ּIh~1Tt^Ev��g�JP�$�|��h��ቇFo'O+�9	X����O(.��S5�n�m[�����z$)=�]�db���<
��<0`�_sѥ��2.�t&#����w[�h^ޡL��񍳨᳁�m��q�)�����[��K��Ѓ����v���?1���ԞՖ�O;�'�k���Ms�<ȹF�/�:dV��~,-��j��D���ov����M��Jx*{����������:Y�(pm�	�Ej8�"U�w�U5�vb�<*Xc��s@zy`);���g�ޗbq��iȶK#�cJo֨������_p�p��%C��50��#��-7:�kOXx���-ɐ'����5���U��кϨɾ�v`EBP��J
\��ɞƳFZ���IJ	OC-����#f;	ه���i�|%���G0s�]-J%4�3���\��C[�D3H���NDGG<�"��Co>�/U�1"���^Cy"�c�Wd�o�M�@�}�Y:tH1L� O�b#�扺���1�3�M�an6��}���-� tI?Z��%���)ϝ
���
V��s�!|�=�_y�����A�.�`4Lnc�Fc\w}fG�`���Y%9���{"߶��>q�6`��e�X�%' ��U�ް�	�< ����1d�W�J���3}���gՍ��0�w�l(�X�!�ӗ7���:3�����'����>![�vf�>��q���1g��6t�ea5rUr� g\�m�W�+#��=PE�`M��j�i�߷vp3�{-d_��S�gW�/" �����#��"WGڂ��L�Lhl_@��f&X�)�Ά`K���,��1���~���b��0��:8vU�Z�͕�P��"i�v�P��GP�}v�#�1iK��*GQ:2��0q�2�(��S)e���p&v�O}g�m�́cM��?��=ۻ�O��a� ����ƺ]<cW�J��[`Y�n,�n�9"���\<A4A��
&A��ؠ��T��ٰ^s@�Տ�Q#.��-���z�ً"ڌ
*^�	ބ����W������=ј�~p��Uɹ;�|C��a�!w��h@�9:_2M|�Ry5�wɗ�������2 �zڧ3 w��G���p��cA��	&=�˪�a�0�gKN�~"wQ��EPiEKo��3m)�<'v
a�h���D����L-H�z��]r�z�j{t��-��1\k>���m(e�k~7��1[�����)r����K<���t�-~Jj"������I�K����z�J~��c�<�� `�'v�W�����T�Ć��U�w#��9:��c����5O
�'�x!��US���P�4WR�5T�E@� �� 3�x���)�(U�a�0~��S
��#��#EO;�4T �B�w����gº|q�d��w1��tsS�}�`�I� 4��>nX�n\^ֻ+ � �c���z��L���3��#�LMES{z^v�ٲ"ň�����7W8KkF[(Jl�+�f�8r������t�6-������6�+w�R��������V�=>����rF9� �S�*�!�O�cT��C���)��{T\�39!��3��MN����Q����r�3�i�� Qd����(�~�|$�$��m���Qa��d ���9{�투�����g��-��Y�B��{:�>����Q�$͒'$J��g�jJY9�[���W�I���@K�xݱ����]�+��r�1��PS!��/�6�zXGl�9�R�2��X?�����8/��������/Î7�D�Kbu��>B��������C�#��K6��9m6d���_9(�-:�<���CÛV�߹zBD�D��J$�<��M�v���h�hd�H�9�u�^�T��"d�L��%y�.Z�~�kD�_�`�4�ܹ"��`EQ���YЁ:�ULQCZ#\���f}�,�F���b�e�TԵ�������`:�@���&=�KM��l�����}�`#<�^0]i���I(^]2��[~������es[jR�yS +`C:v�]��O�	 b�LR��Z��֨��[�6�D��l�?����Q(��rW��e'��t�r����ߣ�kp�M�y�L=�	B]?�^�]u�-�;P3`p���K(7�E�c}����<4��<�U�L6��6�Ŕ48�5�_Y�F���TX�@�|4�n$���
@����M��D��d���bf,V�z��:��ض�hCop-F��d!����fD����� _�i��`;
����k�b�V䦍<���Vn����~t�$��9!�c�]q�+b��=3�}�8��U(���ji�>΃8�Q�mI�6ߝg�CrB�d�a7=�\���+UX��p܋ݭY`-�ռ}3�O�dN���(@"�B�X�$�)ę�.u��r�=\�'��q�ah���3�B�P��HF�Tʩc?��Fvl�l�,h�A��!W��g�ӽ�~/		�MS� -] ����d���Bd�b��@_����>��� ����ӏ��� s��U c�Q��[LΒ��%�(��b�K�$%Ɖ<�6��M�(��
h��dpJh�x�ՠ���A���]ڽ�/�g��b�u<z�N�]�գ,��H��8��HĎ���D�	�� ���-���X,����d�n��]`l����P!��pgrNQع���NP���/���l� �].�f����T�%@%��3�OW��kn5��-ؾ�
3��TOeD>�Tl�u�7o�T�aW�X��>y/8��S�����q�z$V������Pq��ϣ�"����\t:�Q#s�ڲ����������W?�@I����M�|� 8w��|�q$�Y�!�h.$EB>�����G�Px`\S�g�{&�+�S���-q�߻BJ�O�	׃����"~��ͬ������m���k�X�����g��%���_����ntx��ea�K�SA���M�:~�*;�;n�[�lK�[bs�����_�aɮq'`*8�zv�o�k���H�̡p3Q��.M�;=��M��P5�����OxaSJ/wB���0����dRK����T�x�9lz,�#�Z�֧5z�O���J�6�U�Z�;�-r=�q��~��43>o~%u�<0�/6��ZI���X.^A���L�����LY�奮�"��~Z�"A�uU܊Ր#i�W>��#c# �V��R֤0V��'O2h��^�z�E�E�d&�Odlv�x�@E6�����ݕI�����Rkl9�y�_�	2���>d��NF�x[��-����E~X
=�`�vnfv6�����-���DfM���	�]��p�����]Lǉ}�>����3@��w���c�U&5�s���؍�b�!I*s��$�]��"��b��1�cud@ǰ�I��"̮D�ڢ8p�c'�K@��-��Qm5Y�������'W���M��
pC��,{�����s~aw���R����@I�h���%���Ql�a�d���Ig�����G�T�W����7sp�����������
����d^�cK�%M����^����4�"D �ν�����s�S
-���I�l��5�$�g��V��|��u=��Xpv C������bF(�n{Z[��/"i�{XqoE&��X4#BUSG�_����Kg��4j����K$#�{'g|�)������%�Rd$�.�4F|_Z<`w�@��b��IY�A�Q��!�܄+!Z��,V~/Ը�)�4���z]i�f���}���%hU������Da�������,#��q�{nd��gz�P�|D��0V�#�U	#V� ���G)?���S�:ћ��S�Ѧ�����v�K���x��,��5�Ā�e[ +����zv�lYM��Y����"�Z��	l���NsF�˅� K���K4��� �,�wfh�nCoy��H��I��仨âV�8z��ơ�[�+I�܄�|*���ۓƣ���E���6R�^౓tH�*���W@i� �׿S�}� /���YG�����ԘfZ� In��ER����A���
c�Ũw�]�ai�r2���ў�X�������%h�8����У��T�xE�S���O3[,�˱�'�`�E5	�M�}�=ݱ`�n.���a��:�ܳŀDc-��@�N�1�	��N�7""��\{�k>�$����)g��d��f��=��OzA����P�lY����4:C��;+r����V���-?�S�>*C���H2:D��-��#_��ʣ�H׷��\5�Gx,��->-���m�,��!�P��Wj���VX��V)�Z�]�_\u�z�t�G��g�i�`�zߨ�0ܞ��v� 	��q�'�1$*�ؔҨ���養�Dtķ� �K͢���<4*���&u�g��.���u�ʴ6�(������R�1>��~��.�Æ�X�0.̓��ZD�]J��^V<z+Q�'���"XwlfZ��{J����?�H�i��;zm��x˺ �[�n���*��@E��/R87��uWgP>z�g>Մ	�\��i�YI'��^AėrT{$��T�c�o�ޛ������)�r�h�
�oGz?B�-R�+��Ru�И|��v*�NO�#�t���+��+Ē�n��$٠���y1��NLe%�.�u��tQ�oW�F�<2�V��F��'�#��- ��i��l�*r�Py������׀^ ������hr�%��[�j��O�8���n�s���F�:��� ^"�hǂJ��hX��<��Ց�Ii<�n"����#G���BI��3X�[��g&n'Ј ��}��ĵ��*�M-#�pC��OH�o��y��s���� dw��2`�Q;;5O�,�� �'�1p��E�cff�@�����>Q�{�B��f��0�WX�&�f�/�7l4>֑v�=� YCj��;�ܥ v���{��mÅ�{�<��i��cR�܌�a�����K?�Ľ�����o<U�5U\���Y�fCU6Iu�ÿ�	�lL|j�h,��3�ף��.Z���?K׷����
�N���[���w��Z7�w�\��٫��Pb�0��k��0H��3�jJP��kv��,�7�'�V�e�&��H�ӌ\8�>�}h��*��6tj|E�����JZ� ����/� ��)yf�/�9�B�9��_���qGrQK�Yt�I�=ªtK�����_0�q�G�_Ͳ_������ΫpӍuoC����+��5�
~3����ro�>l�]���*����ъB*�і��T"-���a����{rs9E������/pb����Ѿi���;c��;� �|MZ��I��9��LN��8�K����gC�¹�iz�5,eTҔ�,���
G�f�P@�jwnЋ��Ǹ�9�)<Wb�>B>�LE_��;��ҧ2ζy���ܕ�� �9:g�ΘJh[��D�F[!����r3�'�5���X z�,3{�2o����-��ǆa8�?�ܕK0_.m}�z�Z�I��Y���`)�����P`(Q��L?d�NJl��Ĺy��Gyf��V�����@�q��g���?���l�o�dϧ�n�ւ:91u�1�Dz�i΄K��I��X
�+JQ"ק͚ߩ!�9j����Վi��zr5$ש���>P��Wl��X��Jj�?��y����;�3���ˁ+�ق�w��c���bZp�PU���M"���\����(ȶ44�K�T��&k|�Ű�5FĐ�|L�nT��Ԣ�HnrzU�4��[cfe�lA�t~����tA;7Rf��e��J�I���e��yHQp���f�V; E�`�^.J���vd$�M.����!ֵ�<�Ux�@]�h0��Og�� =��׋r2����§Q��ŕ'�ď���,J�9�=V�OME�QDF�vA��j����j��z`=<a{�C�a�}G�r�7vS�Y�_��<�w��0'/��L��JSsLR���2�qbu5���� `���d�ّ�^�J(�	�3NJ����A�j��e]N�y`e�&��ꩾ�����C*|����aI���M����u{"|�j=A�˒��f����;��Q����~�(���&�EU`F������-g���_����_Ma��
�7b�G�e̙�]��:x�nPoG�]�!EAy�Hȷr�גV����/���A���� �q��ӟ�:V�tf��� 4�OZ[U�|�h'E8��KDl׾��D�E��"5��=��-+�kp��潦���/46�_��w]]o�B���h-������¨[	���4И�-~�O�;�{%b���s�ǉ�y����ǭ�aP/L}W�])�"jZm8D�+eS^�0�,g��o�u4��6�Se�g5�OP�rN��<��f����F	�u�V��ÔE�������V�e�p5+C�O�u�p�Q�2H5j�I��mV��R�Cіs�gϽ���[#yz����]x��}�b&t#�;N�nt~��+����c��!��:�!�a5CƆ��Dn+�e�_�.�/D\��r{VD����/#]{���ˀ�( (Zgco�k����lL�R�+f��.�����Z'$��r�t�i��f��%XJ�f�*���}?���QB|(�0{TW���ZW�O�$��-���K��7�dM�N�;:��v)O%�zQ�O�s����`N�|����y��-�ɐT���{W�1|�$i�������R����禈�&k�;�ň�|bM��1��-��%hZ�qU�k��"��k���3g�ss�
��Z�}!4�[q({Q�E��f��o���{#��B�t���"#KO����az�	L�s����v����"�w�NWYF/ޔ����F5�)�;+T;�7�k��F���uv�M}��.��E���+~���/gN$A����P7u�`(�͒�P9���kY�����h��r�_\X��A�E	�����F���k7�)`��0�C��R�|=��}�ct�cHmvZLz���$bJ���侫Qs�`G^�) �k`%Q�P,�4`[�*��i��e��2
��\��9|8i	���]�,���T��Q�.O�(ڼD}+̱�"�w���bV��N��9�Ԓ돲�ŰQ�d��hX�h��{2�*��d�^wU@H�}d �x"s�L냨���>-���~����x*�%��W�����p�	����C��������C{�g�9�����$l�����9���E�=o�����9^쨉�5�ij�3X(��u�1��q(4A�<Q���kT�.u��`'�w9���K�;��ie�����w�q���tKxB�fuM�<��M�H��y�d,̳��}d��MY<�{t��7;�<\6��6����(����aK퍐��X,.�A��t�J����gV뉛��Oˣ�1����T(o����L�.G�kH�Iʣ�۫���TP�>O	����
���h�ʀy�q�x������p)��R�?�5�G�{��Q\��-����+�%���jpd� �^Y����F7�����V��ge�t4m¢%�UYz���x�T���
�k�ub�Q�D Q�
"4%�P�"H ���'o�ں(5*5�G1��(�qϹ�H[9q���3[\զ8)0����n�
��n�v�zN��:�]ݐd���QU_��.P1U���2v�����a�V	��X��ǲ
��zl�3'[&�K!�W���A}���s��i�}����� T�V���)�fC(z��ö"tߛ�
�2�&��(��̸��ME��X�?V�-�P�Eb����$|G�tW#5/��v�uAB  ���E����*�QWCw���*��`~��2��j�AyT�}�3��S��H��u�W�V�o'"�=UE���Q1zKj3������oFE�,�޵�I^�#���k�e�����|�
%�,�~]��sln˗Q�hX��L�bY"� 8�ZŀNܝ���I�\%E���I\*�Mi�V%�e��
Ӄ����z/�	I� K��"��)��03��mcZl!�끵����j���B�8T�t���R��j���9<Y�2���E!��n�$�RBJ�<���nS�*0+����xf�j� �:<��W�RR�{���� ��3Zv���Ut���/�t��kk�8/E��F���B/Ab�hJ�g��oӛ��ؔ���Ee�c|(����NP�5�����C�.K�|�Z���e�zj�`��tT��O$�-��!�q{n�N�-�]�]�%�>9g�����hl�*N���WT��{s��D&���qtaW�Jp{���o�0����{�4u�W6$Q�+́��d ���k�Rz=>��̥���� `_�ȡ��E:�7���wn?}�X~�~Ϭ�����H.,��O��ey=\)���*>�lC�����ʩ@�4���W^Q��Wq�d��9����9)�	>�<R���c�����B��?j��g.�M��/ԇ�45�Sʶ9�8%��Xח�Nȣ�T.�&�v�l��3?�y�l{�b�m��Қ
�'<��41���l3Cۨ8�ʪ(L{����KOLc����d�H[�?1� �=�}��!�| s��9���y<�o)N���a��	��t�`��A�le�U�f��ҳ�7���`�C�!�;r\�V�&�FRȎ>$�.�(J�[ �0�y&�6�R�S=*�G�m4�z)e�q�ͻի�4*��T1�2'�FE{�klGZ� ��;���=s��0�PQ7����D:v(�#{ǔ�Ư��7,q}������J|���ȣ������?b|�<���͘=C�<��5v��x+:	e5I�.Վs�G���)T��{ ����(NT����� �;e���|$�ߖ��?���>���0�S� ���r���dn�P�*/p�[�/���auY���à,k�l5.�ֆ�zQZS^�m��kK}`�kJ�WSJ�n�=ނ�a��y�I%"������#�Zǋ��7W�
+�3ɒ�>�I޲^a�9z����~ ����	�(cjL"ہ�9Toʮ���B�dT�+tN0�����C�!�#Q��Lz��'�� QƷ/C�0"���aWVp��.���"o������9��������א���T��}i�W7�9�jcV��8������/.���jNG6#4�}K�0K-���C_բNq	u�>AW3��{h���Aj�0>f���+�o܃ ף�E�"�q��ŝ=� bE?��b���O<[�xb\�K��6�<�"PT�bȐ��?im�9�Aʟ��0H�0���+�'w��Y��#��Ol�b��y
��6a���i��C���=�����b�=ۺ����PLK*%����=�k��W{�P�l5T�촞�
�w|:F�a�rĀ�=������4�ӂPF5�~\���aI�&p��7(�����C5�2Q�Qe��F���~Ƴ�� D=��큠�-���|3�e�T~IN��Mf�L�n�0yơ�'>m��'�RdF��#E����s�S�T�!L�L��/�) �d9ȱ��`��2�t/���2DM*���Hv��
�^�-VbL�k�u���o��5Z�@�R��ـL�(�Z�̲%<���ٲ(�OBH�����bp3��B@ ��tFX�#w��&
o37�}��L�J$��H5�� Æ;\��.QV�IY��#:8�t�L�(��gzB<o%�!�;��3W��/�ER�7�X9��uߋm��Ƨ}�#)�

"i�@� �?�|ǅ:C)���&s�}��%ق�սX���5��셙~��~��Ύ�h�G0ct�.��C�^�r��7M'�_uL�˭2�4ΠS�,!3�FL��g���.� ���[Ǉ��V��Nܔ7���/K|��P��E�f�;;t����V��R����ꂝ�@'�Bm
;�+���x_m�y�]HBe���Q��S����Q �B��q��.^�N��$K�pG>����{�W�Gs�J9��غ��}�y(�p���P��PIKβ_0�A�S�H5z�qEk�E�3÷(rR�_�h��i���H+�NH�c�C��W]����Od�7/MZ�3�lz�s/��~Qk?�wIr�5�,V��W ����] d�T�t��=R�m>��fY�*�	� єC_���c=.^����Ђf���a�ʹ��8gqKp���#�q$+R�<���*�@���u)��Yĭ9{�,��JKpL��:���' W���M<�hR���b��M�55Z�9�:�H�1���~:ȹ���G
 �:�'��!��j��~�(��h�R`��: ���Sv[���E�y�:l����:m{H���:�ء�bͰP9��.�F�K�5�Ʊ�a��G��sC���6+,2��,�z
z_F��/Ah�=(w�H4�P}��y
@������-��O��)��N�PX��1eE>ް^t �_7�X�6��h�4�����A�cӞ�$Yz�[1(��	0~�C2��y~VI�ӟR��D3�����\z"�٦f�u_��:�����0}�Ǯ��)���A�h�5�qs�΂s>����(}��j��贙�_Y)�;���uk�}.��o5
��7/�-$f�=�2���M�8d��B�@��r��=�E#:��)5F���%�}���#�D���^�dOF9%$.�22Ѐ�m-U���Z;>z�:֕��c
����9FZ��Ծ]����mK�h����K�i�f�etUx���׏(��W����o4
f�,��q�7�[�k'���8��ʮ)=ɋ%�n/�z<�-�_U1�����x%��hT�O�k�`� �$�D�� ;_4f�tuOK��݉���o+��$�}��в���ZTK"t�KL �����[Ni���r3�N"*ɒ�u�N�TR[N�6�v!�h�f�;�'��w�+T>�'��$W�z��[*��V=�j�t�\��U��s\���Q5H�5��� ����������A���g�V(�t烠Nd�\t�=�Çl��n^����L�n#��50_�ʉN��db��4�r���~&C;N�K�J�Ŋx[���W�Q��ְ��"^�Z����O�� d�^tFŭ������n���$D��p�Z��`�4�JOY�s��`�=�A�j�>RF7���^�4��쨸k��t+��-�r�3#ݞ�>=�����9<��51'!	W]��ـi����X���બ1=z�#e�r��x,� ˰1�{!����p�b�� ��!*I^��.�j� �x(���<U_+�R?%�Cǣozh�;�'�_�<I��Y�i}�܀PHn��?쏨HϤX&q��[��|�=�0?<V�;�G�W�'�d��B���h�z��h���8{�ߺ$b�J�R'� m�[�,���,�S��H^�
��<Ż�g9��&�� ������"y�z����I���W������S�e*�iT��ô�r~o�����m�`F�O8��; �����Kt��3�>��tx���y��2Fo�{9�f�(�U�ɘ��3�T�����ô���&�WdW#��������4�ުd�MSp��pbY�qv��{N�U�P�caKa売�e��-s��Ӑh�bD]�?t4YZQ��N�g���<^]����� 	\�K���rW{<�^K_˻B�@Y�;P�sh�-v��[T�b/2���T)����?�*���S�� ��VV"4�czRH���ȧ���"��p��]�.�5��e^Y΍HN?o]$��M���=gȄ�~����]�_�~����?~߄�{BOH؍��{��?�����[Xm���1�	�T$��|�"���YD֢!�%���L�o�dG����#���ӯ,׏��Y�;����5�I7�:lR1���ӬŮ��.�'���&Ο��~�[�Q����,�c��~�ي�O��$iߘlVEtk~�@TT,�1��\hļS1+.7�6���~z��1\�v**�P�,A�!�=˧Gn}�?�9�=�*�}m��N�.����s��C�H������S��3��q��R��h��w���b1)�#���~�c�zX�no5n�}��qȓr�
���Q�}��sK�v�e��Ro[+��:X��3�3E��F�M]�O8�x�����dl�S���t ��!�?�d�H�#�zb<OhYoǮ���.�qPf�ٹ$�i�T��IPS%��0$���\-��^�܋:[�$����>ҁ��'�~"@+nGrHu9��A*<�t��O]�;���P�2�-3����_�#'i�m�Շs��i��W�Ծ_��>��g����ˊ�~�1vll\`��0�̶�n�:������uO*�Z�F�>�vH�?��2��$ƃ=s�^[���UK��T�4ݞz��"��y�R��գ�n��tO4Q�N���l�B1h�o`��!l�ad���oX#��\��ޠ&ْ��`j��˦�.rU���Qjo@L�L����ob7r;҇��-�u�K�����I9h�xGr�����c������M�SN��
|�3�U}nO�,��?��ߔ����߱�n��<�Ai�2>!�1�1�@J��D%�����HYҾ�ެ&?ΫH�Uі�8��T�m�	��q>3|���qFU����S�21��r�ۂ}_�(����C͜/�TpAV��L��}rD�Te�%w�d�BYոq�[���0[z�o,�7��!7�)*�ܗ��X�S���m�G���;�t�HC��?w>b������07C:��@�کj�k7����� <�\���)��.���tx57V:�6�h7�hz��'��(2#b��W}~0�0�5�:��<�.߸�
k�u�8~�>��1Z�epO����v����~T-��/[��U�5Y+�Q�Y����Xm;8U�ݺD��O`��Z�����<�CE��+�g�o��Q��h�H��I1X�(�>
�Hz��ʕ���ϓ��� ȓ�e���J�(9A��)�'�hx���R��7_����5C�ɂ�v��{S����li��)��옉Y��)3�RP�[q\��h�Rw���Ӝ������LW���%U8:�?>Ж@.�ț�>t2�jk�m�#�d�y1氞�E���H��X?�Ţs����l)T���X�n#V�#X/�]Zo/|�/�E�_������BC۴�%"d�<��f!3v�Q<�Ŏ-`wd	x՛�Ϯ�j�f~��.�� Qg�sйQ��fb�RCEF���i�ѷ;Ņ�Q��$��$\�'�g�s���,��O�W��f,�a�~�����'Ctϯ�Ed���s��x<��ꪒ�a|h���+��%��_�f����	�5%����U�C��j�����f�6x`��!I26��`�K`{��3�H�P���z^:)�@���@i��{z0EF[2Ob������C��j�Ku�4tXJ��*J�&x(�>t)�@XC����ogP�$�9�^�A��׷is� ��J���[^��K���2�U�Uo�.�,���[������)B�x����Y��J�E��!����CѠq�'��5�:���	HA{1�԰��w���%K� �˄j?�_c胋��e�$)1X_�ͬR�ײ�zY�c��5�ky(.�Ay�7�]|���F�FU�P'^)\k�Jm��=m���\���?iT�@DId����I�:δ=W:�s��T�s��� I�+_R�I?u����w��]�t["��g�,ncȦc0�.Jo���!:�������Bl[Π[W�G$��W)�#��Y��>G��8n��_Ϝr#���ѩ9IV<�C�רn����YXϛ�ʩ�Td,f��H=����-���e�K�&�A�n@��p��xr ���w*�3W����kj�U�),̖�8�2-�SRۍ��Մ0S��!SyC��Ch�"{۾^��Y��9yݭ����!��m��D]�{��߫��j0;����I�&�������F\!����!}�0����9�X�ô�[,Il�u.���=@��j�� ���C@*�MM 1:qP�w|�ӫT7u,k%pיU�A'�M�W�w
B�}��i��#��
���"�@5�N�6�xD��H�)4Щ����9`�5ĥ���ӂ\�j�F�8w<��2�?G�W[����o�+��M��4�k��x�v���W�a�	Юߣ�F�����Ԭ�L��^Ty�W;���r'|Y��o�e��i�3G��-�H��<��ýN��Cqk�ps��%��q���:���*[YL.ܤȕ��FB��R�)(^����Z�DB������M^����G�1�Oi�]mvM�Zm֍7{p���o��I��R��'Y�ķd�3������&�a������x��ov'���Aլ��k.|`i��趘/C��`~6#,l�+��>ۻW��y�� (b�3f�С��o�{�v�n�� ��9Lo��	p��,��%[��Ɠs�\nG¼�LEr>���d��n@����js�rS�A�tp��
���3ou�L��?d��R|�ȃ��Hmq3�B43l	�#��B�@K/	a��tL�37LMn"�th'F���3�u�b��R®e�r�CvT�~���s�U������{>�]�H`���I�R�-�W�(�1Hg}�~��u��I�
�T&<�����5L���n$�H��hU~�G�;�6��!P6'�k6���1�,�l.`4� L��B:��W{h�
�����͸	F�.�q��vN��T�?�TŽ���{nf������]pw�����֙Ϥ��-��O~6:�yȸ!�m�ςˉn�"�?h&I�ďy���&P���<�]"vP�}���a�L�i� �W����6��n0�!��ܶ���߅�hg�9Q�/�2��e|������(�[��Ld���,܁�Z�Β��C*2�u��#X���QK	YI"�����]����e#���� ������d � �5�[
���<Y�]�J�mvr;���{Į�T��0� o��sϸ�@1c���e�����>v�'A�&^a��� (2�ע��&щST�^�m�!��L��aw>�?!��3�޶���ў�����_OH���*Q��,�о�W�'Xo�n �?K0R�3ARӴ���r� �����7��j���/�/�!��V$dE��eU*"��]��`��ﶖ}�:M�3lե��]�2qydA�l�=%���15+-�z'ޅ*g5�L�No޾��eܳS��g����^a������;�o}
�ٱ���N�&���O��;�{o M+u���G��ƌ�RXUY��������%��� �J�����";e�ƥ����*�3k�"��QU�_l����ǐY.	���G�Ϧ���`sy��e��)����������ʙ_�I@�����"�f,�a5k���LYވiV9��i_���]l�kYt|#��U��ҀPP.��I�dc$�����_�h����ԡ���/�@e���A�6��B~�%A� ��>) B'M��ʨcˮ4Wq.�-�`�<�'�b-L��P�?���y7zQ	pgN���_��_���0#�fS�{�%����<b�,����M��`�N��(Q��)6Hfy�N��#㈝�~/���	Ĕ��*>��$��=׷��7R�ul�Y������
�8�p�3��J _��G�L-5m���_@���"	�C�FGz!�MM�`�%�f�Os��=�z,���"�)
m�a��Cqm�m����*P�\	��@��m��P��\�]�����V@��E��pw�y��9,���r�--E�A���yz�Y:��V������/�re:��N}k�����a�h�)M�@X�[���:�a��k���+��ՙ�<̫zf��K��������Kr3���N3�G�UU纀$��%X�(yb*MƲ���>���ۦL�p/��9��ܤp�Ԋ=��g�;�*Pi� u D"����%����w�*�BP�Z9O>�+�i����z6p�o�i`��,\������:�n� ���O�Ngk* յYku�I[Di��S���Ǭ��(�1Y-p�+Rv�ij̎����׸v=��ۂ1y����f�&w"I�{�g�ؤԡNp���{��Lt��XG#5��i8��b��ȍp,a����\�ZΔ�,���kƂH� r�x}�y1�1���MU�~���g��¯W��`��#�!�z�`�:~ �UV�zA"`���xg��<֭6֩�US�i�c�J%�|@S
?Sr�Xzq��*CF�U��)_�=��Z�S����\��9]6M1��T�С5�s��=���ݏ��%��R,��8mk�!�����aJ���I�����Q��yrw�����M蛎���b����O��ƽ-u0U���'��J��d��֟�����x��7��*j��h���lĴ�a�2�&n
��eG1���s=E=>&�����%U�"8��L��*?N-�ɘ�y����8s�XO	H��`����"wT�f[�Rm<�b̠�տ��֔/:<���z|�M��.� �"���n��&aV'8�,�/�M-�U������Y���t�2 ���ȜUt�\��&��3�s�2�����>LfTlf�S�GoQ�O����go�\j����O������_��g�y1R��F���i�� �#�F������D�Qz�"�-�`�E�w�#0hE����9zi+����&��҅~�S���S5!�	� ��d�GY7�﹢;�-4Rb����8w����r_I���N�ʠ,�T�Gl]�7ʦ���Qܵ�-�Ʈ�u0a
Ny)L��G���|�e� �#�78C;�BPM�\�d����h�x�}xe���Ѥ���9�;o��o]���f��|�Y>�X3C�� �|�����r���)�\ �.^�m�lf�~�,7N��B_GJ0�-:�%Q��F	aʘ�y��K�˖֯б�
6^J�'��Kr��ڝ-txq6)1񠶆}ʔ*�*g�}R�L��7���ܺ�{�-���Bb�ds�׾��c�I@f?i�SO�~�$�wtt9v�������b9�GI6�F�"��o�!��}�ªt���筞�6+����A��.��oآ�6\�=�
C'�^{]�Un_�=ږ35��	��V�ڞP+؀��=D�ic#dEE�袉�t����F���')�/x�݉�`�T�_I��'��+�d���(C4���{��ƚ�ؚ����)�؂�c�Z�n�Z�Ձ�ڈ��ÿ'�����x�`�3�<�xX�Ҕݷu�Gz�ķ�������˽X��1˟C�����`��g"<�v�m��<��<$@y�)��dA&��a��2,JAiHIb���c6
&ӽ��v�� 5R�RѲ�I��3Y���2����S��K�oY���N��V6'��i%��X���ḚX�yT%�+�䕏Ȫ���{��^�s��9�ٝ}�gs8�e�T�����g}2��N[w,�#��:��M��������A ����9/��� �ǂ`�w��jf@��J��js���6��� l5���i0a�����Z�׽|`�UC�'�Ye.���"�\v٬���!�r5E׿F*݉%S�6	�IT���Ifs�z;�=a"D 7��5�yZ��17 4g��--*W|dx��B,����,S�g%��DG����E�������+ai )�%J/H�sC��IQ��Z��AF����j����X�͖��kߧ�<=a�	qi�:;K��*�4q44n���{�{�=֚�n��6:;߱2	�����t7��|��o�����.���8d��f��mg��]N�����)@�l�&=IG� 5�W�&�,��P18m��2�Ǝu��<�$�T������[|,X㌹��<ԓ��y��Q>@)KS�ѹ�+\�`�:S�-��	^�n��V�	7�>x��a�%?�X�i��I(+�.T��7�	"sz���EO������؞��"^�ٲ�qc4�n��y4Eg?�lPAr�8� �w���~�<�&��u1)'�)�'�z�=-��F�w��ǩ���糟'�Q��QucUԤ��%2DO9br��(6٘U��<�Vj��N���}���I��+ý�H#�G9������	Ze�w����Q��K�O�cx�C��m���FJ�v����4ȖD�?<F��pG�h��۰c��.�)��|���T!�&��������f�c��#�G�yJ�\y�����$0鮦���l#8�s`jm����įޏUuM�W'��|ۑ��i�
��G&��ʪ��;ݫ=���5��yo/i�~k�~/���V��F�x��N�_��ˊxRY#:�D����N'�{�v�]�����b�P��W7��~n�C]K�|h/�5�v
1�j�SsMjt[�T�{GÊ�d��K�R#l̎�	Ty��ue��zL�@�S �*vgT�u����I|�
�$ZP����-ś-.���[L�#��|T�-O1W���b�A�fI�G)RI�Z���i	l�<��tߍ�\F�I�8��?g� ����+�u�m�x�}&U���I�9~���>�Ք41����D�m���T�.笳����g��tf���@w�E=��<wh�<76�]X���2q[����%�U�-{ҤٚP���,^)ܧ��$�Ф�m����[���z7T�������'���bN��qC�0d��\T�6��2������`�/�F�J�q��.X��r̈́0�X/P=L8�۫J�IW��8�ai|����BY��!(_�ظf@T��[&��;.e��iҐO}F?��!����B��1��O/9�K�_Ҿ?[���=	 �p��1d���:��؟#��e�C��W'�,� �i��7�}1N#����w�L��!�+^e߫D�O���wL���%]���}�"��cg*bE�EM�%tڌ���o�-#0��[Z��7F��c��������PɆ���Z�:M�E�A������rٻ��7��Ȉ��XO-[��z4��u쪭ᴰ�ozԛzK���w������Hc����]�^��`��gĪ+_[�4��.�)ͭ1\����y�.ԫ]�a�8B��Ӂ�|�^�X�{q�1=P�;t�'HA�# ��A)�;�i��O<L�ѐ���ϯ�K�$��S�C�%eh�a?]N�`5|��H7�@KD�R���͋��A��?W�+����U�iDЉ�����{dӜ�D�ET����yQ`Y�<Q_�������6��E�w�\'�\�L9�f����w^*��*��H5/�kXƽ�i�� �g*O�/�{>J	@N>��� �^�����rD�Zt*�v�D�t����!�}�eӸ�`��&�NhV6u�ʙm�Ѝ�4:l���oW�Z���c�4l#;l��&�*e���\�YCy���8����rlc���AϣD,�߯{�Đ�w�o���1�]Q���c��T#|�u1�mo��hi��R��f��<l� �Ygd�T� �EaW�־-�
ׄ0�,e���F�(� �(x�j>��BM�D�
R�܅�k���>A��B�~�~����g%a�50��N��q'�},(Q1r�o���_����"�Q��/a����c���k>N�tp����
U���SvX�VG��@�	5#��ya~���R��;VR����"56T͉�?���lt���@�<ƍҳ]r����1�-�L���l���� �`������/Xݹ�ڻ��ā��"T�T_S�N_+�US���fDv6���SG	Չ=C�o��͆�6/D��O)��xXB�`5�;��,�eB'>��9����>ũ�4|Mj"�V�\Chz_�3��{\M�z�:�=�o.�%�$��j��+���i�BH�a��Lg���{�rx�W�;�����O�Q����~�|�8M�Nl�VZ����|�Z��d���O_�`u�V�h`��v�~Pl�>o�W3��~��F.$iK�<�sV����Yu��w.�ﵰ�ف��VI6�=&���6h�0)U�"�.����� m�Y�S��v�RGY��0Eȹ&� ��6g�v`����-��D�!cB�ӡ���x4�x^\�f	Ym�?��&\N��7>���ں��6~��������B���On>�Rn��e�e~���i+�{e?�N������NO�6�"a���A��8�2O���Y��S��^Ŷ����zw�H:�zBtl|b���f��B����Ök@СT,����{eZ.�n�yTu6n�	}����y\�����\��og�r��6�/��J4�NJ���YX��(�k&\���l^_ӗ�p�ls*^*Z��WiˍI����2{��"��X��T�S<�0?Y��d�/���s�K�&6ɩ��|(�Ai������7��(u�U
E��,�� emd���%�"\z���918�7�$�k�k�Ks���rl��{��'����EZ�RS:��E�F�،�&��t,�a���]W�f��$�A1!]�$��xdA�Vy"1��̈́A7p����1m���Q�$�g&�p*��B��������jf��۸.���bJ���JC�T�/K��_�F���CY�޻5N{ZFnV-_�k�>"��Uz"'o�����y# G�j$5���
%�=o�]M˖��lR�cNv�,��d���8�� <�u��^��S�ۊ��Q���0�$->ڈ��馢W��-�Π����Ԩy�%�q�@y�|C�H~>��(?+�P̌D�|7� ���&�U�@�
0�Fx}�[X��F2V��(|;�6���"�T��eL��ʺMdc4��p[���:	T�N?P�I��~�e�u�&U}�в�0ɽ_HXv�8���%�p��t_'���\����*>��ϗ��Y��D��U �v'��mr���'Ԃ�8����fc�%���[��BǄ����1�)���	:��J�@ s0ت�b.��IA��8��������o}��$E�6�4�|Z�a� ��'�֪�Gt���B�X�P� +f`��׳�F#S��Ee������]��"��R@6��6���W1}��Q����L��(?�:��7Q+Q��S�X_�_� �s	�"ɐ�"|���1|{[5��oE[��������g�|�m;29��hsT����Y�[غI�̠=��BS��)��_�9���-���=y�T*��a:�E�O.8�U{7�2!V����{�L�Պ"M��^�^(+��v95ͤ���c�C��a����

��l�@��,���,��"�Ĉ5z���6��Jh�aZQc�B��($�&�z�HbA�� ���ݨ�{�]^�֮�{U�'V�b���i���q�6w����R��\e��l�~�*�6,�͙��s�/��pO.����TQY^��*5X����O,`N%S f�厅��)�bF�B�
�u��[��U@�`���8ՆCgM�.�N�۠sw�*�a��O᫡~#aeNcN��{_ ���*�}�
*��tw�]3r�y�}�q���i���ś<!}����o��A1���'��W����n彽.��ð�%O��s��9���]�m�89���aXO�g٭��E*c�-����G����DO#/��n��L\\#uΌ�*u�7RQ�Ĭ$4/��rC��jҥ���j� �u��wсX?-|�p�=ټ:�>��K��҃^�R,�W��<�֛��w����R��t�Qmq��ۡo��� �*�(��k�ԋ~�&�3x�8yC	Ji�5��‍4 ��9�������k�(��3�g���/Cږ�)z_K��O'�!޲���zC	��f��:g��ޘ�7�4���rs^�HVW�LΞ�n����}dX��T����<�,m���)�b�˰�ij�i���|W�^�n��:Z����P_��%o��A鷲��I�߼aduX@�����]���~.Զa�y)]���zpR�V7��ہ"R-��M��s�:K63��v��F��s���ű�l˃s;.�Y����#� E�a��C�4M�Y��?^(6�7�*R��9���-iz���i�[�up�b��^t ����:]c�!�(���MV�Ǖ����-�<���g��1 �c�T��
�2���Q8[�~!n�G�Ԉ.K�xa�u�Ak#�����RVs ��,�~A<�j�p�_��ԂTr1n�to��43%l�S�������7a���B��g�n�Xe���,�����|���k`��?3?5@3�I�䖟�B�NZv�/Q�*�Ƀ��1ϖX�	O�i9�a�*��6G�����>�Ζ����,cvW�$�ή4;���ʎ�y�����])͞���ԙ�M������4��` f�g��8Jx�V�l�J�n����j(���d�
2����_R̖s��{��=�P}�
^����}�c�+<�R�ù�B�m�i5��Ԇ��Xz�&R���`;�����B��"0X�-�ں��/in���b���ɐn���'�$�����M��u��0�p;���8�B�w!H�dXNc�9���H�¨qI.���2'd�%>�1>'��9g���}J�9�<��	�i�������d��t�և���z�m6Dj������{	u�S�W� ��?�%ϐ����d&�^q(r"�t�	���+k]��U��Q�N�.�g�2� �*0Z� J��?~E;l�#����b ��6��W	�9���ò0ޫ��V��I��sQ�:�%�>�����^ѻ�~�+�~y=�#gY�E��ሆp�+�(���;���cK����/WS1�>,�n6J!����"|_�oڸb�.ˌ\/��|m�i�[��Q�㫸��52���FB���P�@�I�1�����$ޑɧ���
�
������3���l�`5����my�¯�ࢎ�<tU�C��&$X�'s)�}i�X��~��fG�vn�x��L�+K����hm�W&��\��c�F�@�Zk�;&��W]Xר�5��4X����×w~�=��DP���,y�9[U������ⰳ���r���Q��������U�H�����2ao��{��F�9�|e�v,�X���I�ϥ�Ѹ|2 �~..,���	`$HG��@hƔ��=%�x��\�+�Zȡ�ߔ<6'Ia�B������%��������ߔ���o��̏�� ��-�z'�d��j���1�`�d��������+'_HQ!��de�9�3���>����Xc����Ф-�"Dm[�i�>R��(q��h��&�P;mzb�؝s�a�$�,�"������z�FU��D}��U!U`��;��w�G�ـ��@��<�F�C�+v�����XY�95����i!�<���8Z]�3d�'���ļ-}~ �k��|�f��+/r�'\B	D/���䶓�{�Us}�z�8ٶZ��������+(�fZ���b��^���kd�=.�����/���lQa�����d��`�I����v�ȳ�D�P�q�SP��jЄb$�0��zP���0�ԩ4=�O�󷜢�*���`v`���s��w=�u�6,�VOW�Ϛ�����"|o�A��O�EI�`׷��D����lhi�e�#��Ƙ�?���mʺ9unͻ^��|d�>�_�(n����F.����j ���g�;D"�~.�a�U��S/�� \q�_=!�t�!�t�����5F+��G�6�z��� �����(aU��BPa��v箌�`�� 'ͮ0�r�������y�&��<�ĕn*D�<��B�US�3#Z<�:ƧEG9D�n���}�l���#���)�� 㡁8$�n$,����@GV�f�+����%�o�۫�����I]A߱(L5�y��@\�������!�_7۴�й(�/�dm()�_Ÿ -1\Ĉ�
V��h}4L������(9� �[z8?c��= j�@Q��[����rm�k���`�+���5��F�޼���BPy?��x�R8�3��gFs�arml�F��R���{�0��Up,�����P�������
V>�j�i������j4�4$fy��}�Ԛx���[�Q����j���c��r��⿳H��-t7������N7j�%I��R夹�΍�������}�D�	����ͳ���[|�Ґ��Ð$\�L�U�y��������{})��$�^gK�a��R�@Я�qt
�t�C>?��>�����X)��p]S���=A��5�_%S��wN)[�^��.Q�ϻ#7��fW��S�8�_C�ec�����k��
�^1��Ď�]jZ��ss TAr���Qލ$e�1�m%�r��}�-�<�Ņ��|�d�i�d%�('�~�=�MOzJ�7�	9Ak��:��Iyn��z�&kL�$uf.�9�d>8Ӌ"��u�>&w��&�[�E>�y����a揁ξƑ�Fln���ߦ�h�C���5��E� ���4gNF0��H>���6j���Wo�-N���X��.��x�"/:�%¦j�d2l>e�ؖ`�yNM��<���x�3��H�L#�q�b5o�6Z�S����oa��
[*��g�d�Q	���$̍yUs�6g�t.ڀ��?�ڋJJ�$Ҟ��(��ؿn؜�b͢��B{�|�E�1k���L�'�K��!���W er=
�b�qʆЇ�d6�'�w���ؘ�y�Z�e�%/��h��9[�tx�b�b@P(Ӌw�0���V�8� &��K����u����zke.��H(��� �ke��f��e��5-F�cP�vX�skU<�RoDZUg��P�o��I�^K�^:4x�;I��L%�*@�CW6�I4�8��3L������R+�O]Z���p��q����Oq����R̴U	����^& �b|�������,p*���e�\�]šK8��F�-���56+5g"�6�5O��P�R#[_M-m����ӲRc��t��d�ٺjӡ�k�+
��@H�f����L��(45�����t�אy�ގ�� 2�ˑRs�C�"�O�7��� )��S�xҢ���Ҫ^�}���⿐N�2;�즰� i�F��e�,\���kڲ�r�������Π�1�]�0X2��9qc�� ,A"㌯���ݴc�])A觽k~L�I��Ӹi�z�&�Ǖ�殭��������K'3^k&o(ӎH�Oqd�*ۻ�8�	5?�) ��P���4J`A����*��HOt��,��BR��B�%���0?J�p�*TW��_���cu�4S��
Pz��D��z�oV��^dc]��xV���"��S� �s�k��Sx���N&�8AQ��L�!O��'�擴kh��|��:EV�H�ˊ��!�ڔ��i�j6�'9$��X@��<�J�|���^�ѩ~���9(Kv�DDe]G=3�hu���X�� gG��'ҳy�����Ƒ��a!	^_�7T��O�*�j�<�|(��9R����e����VP��}��G�9���Ԓ�L�O{#E��U;�&niN��!x���&H�bo�bܭ��u!��0K�+)�ߎ� +Y��E�.���^_��}ک�a�����y-Gj��/p#���o�}�K�ב,b��`y�1��!:�T��)�R8�����IB��H;��W{�N�ٱ]�	Z��r���#��f�wzX��m�	+���}� �d�å��ـ!�p��&챾�	�}(��'ֹ�챡��K�]�*�W����8��2e@3n���C?�n7[]͕�PJ��_���DQ�l�	��@�* ��!)���Pr�kά_�*�]�E����sL����Ms�]��86�mDl�t�W"�g?���;�@��� ƴ�L�@��K.�d��]����7�
x /՛v��}��Yʚ�5���c�M��u"����)�^W+��:3
�w5��ZFj��N�Z�BF���>Hfy�,���q ��0E����j)�Rz�mw���;�F���,E�Qt�X=% !�`���=�)!m{�Q�k�Ql�gXj���y8�vׁ-���tH)RZ�6�3�g�,��yW��Ø���f��k�f%!~F⎅�~�W�w\��c�:��+�G�Gf�H��D{�;&e�'d������#��3�Iw�\�QY����D��Mhh g��'����Fx�������[�p��z��_�Iu�L��/�}��� g�f���}6���Z�2aj��\�􅬀7����I�<;�؍�;�n��-��5w&�JI�@7�)I�D���E�˽`sG�{��8�4�2x�ʰ-�!�J�u�fg�m��h���V%"��e�%� ]�ʱ���h�����-c�ɜB��0)�hk���n1���7�R���uYԿ
-WֻnZ,.;=�S�M�B��?P�br�p��k�gˤ-:<y�7,�}�]���]�-(6b�N�[.v_'�v���{r��(��;K�##Z��V��Z2@����&����<�qH�^��t"AS�3S=ۤ�*�̢�J{��]yIܺrTM���)��d)�	r�����BL�Vw�i}�|%����b�v��^g�'���<�k�-�|y�^;v�O���ജx�̩�����rHt�P� �c'xZI���v�K�,L�7�r�g�׎E�"���u��Ps������=>�{�y���;A�h�,���I���x���Y��z��r8v�W������6��3���X%�e-����2���nwܵ'���5|������x#f�#�E����gbj+��Z��zi�y��zPf�A�����z��|�sP�����W���w����y�i��!�ɞĴ#�"qS�\+���u��vӒv���O�F�o/��1G)9±T��)�]e⮶�SWQ���D�$�����J�����#��TP&R�0�Nx>���S��_m��zTX�/����/��.(��`���2�~�Š?ˡb	0k�kwU���cXi�E��;�UZG���<�d�\癉��05K\a�}��_�{�9���a3Q�K��&�Bg����e2������C��~S]�."z�o�+p/�E?`���0�ürf>G�i�e�)�O7����1ԓ�}���e]�yI^η�H}Z#��L�U�ef����	�~�sܜ��	���0J�v3c(�v�G���[�z� ��/���N������Jϔp�u ��,ସdK���.����HJ~_�up4>�����7f�p���"�4�fW� "v�G��uF���'�f� ~$���Y��f��
�L7ㄼK����u��skܫ��S*r�����r:r���6dv�o^צ�I:F�0tIO��q��E�-��d }PA+�v���MM�|�j�Y}���Ĵ�xy�f��Y�9�!�ʁ�����\�f9�C��p{+�}��7�͌��^P�T����EP��Ac�����
����}�z5�dc�t�Z�m4�Ҙl�� 
;}�1�^4\���-��j��@�����l�B/b�n��ǅt�
6�:����a���I�n�"��I�tC���Y�R�Ier z�_�`l�]���M�i�01���dW��k��!:���i�K�	�Ĭ�n�M�K|I:���$�[�P����ei�����ה����]	�ɍhN��A�b�,>BKN%��ߐTS��h	��ӆ��RD����%�	�m�~K�Ρ߳��@�M�S�f�&[�ip�n8oҝ�\����8xfjã����$-��.��c�n"��-������)��4�Z۟>J8��Szڳ*�kO8�ӯ����&@4���o)<��9�;$㧾�j���o�ON�P���s�]�U��NE�$Xe"c��4���FTx�	�ĺ)�ԉl��t6��aR��kR�x
�-�{�ҷ{Ҥ&�Co���C_y�4�߅��R�?滢��R��la��p��t㐑��K��
��I��R[d�?hsݘ,��~c����{�퍲Wxn���(l�69��OW����<B�m���x�����ҁ�ljH
(��#Ĵ&}I4��+i�����X�N܅)��ڀ��;��y��\Oc �]�`|e�z�*�m�jG�CzĢ�q���/�+巇�I�ص���Ұ	J\��Y/� s��8��l�D��ֵ�2^��N�QQ�¼�슇��B/�HZ0����I��H6�F�l��q��/���D��o��@�O��e$������@� kt����b�]�ȐT}�h���
���Nm�,A�e��H�d.���|������k�~���S]�� \����?�'�bԛkj�B7+��9�ߕ��'���x��#4m(_tC�b�!hD]���ʶ�~�K_��v��Ć�ߤ1�"H��gN+	����4�,dۗ����,!㒋w���!������XYE&�#Q��0��3��/6��Z��Bgk�?�F!Ѕ�[���T��`,��b���J�Ѵ�åW�^"+^��~����@a��$/�� x��\�ZKM����F�ħ�)��n��r��,�	t��h¥%�* = �+��S(�s��S�4��58H�J��s)N��A�ߏ�Dk�[6Wl��ǳ�� �Ngs|�ւ�f�7��T?�0Y��1ĢU�~�SSn~LW�< 0�v�BmՍ��4I���K?��y����.��w��UC����0�:�y�{���K�\이詝��8+DQh��4����1qi�}&��U-�����XLC�~ƹ�P�p%�r��L���
JH�������������
���Ϥ����?bjt,毾��=up�
Y[HZ'W)}��/F?�FZ~����p'�s�|��$�)r���^V�[��<�R2qz3_�2�b�d�y�z��U���Ȟ���.��y�}���l6��T����<ѡg7h�<i�RýW�ё��O�n���n�/��f�l9)��GA	I�;1砀�����v��{���������G�[!�H�U�?Oq�s��v��wࣥ������Ց�3��.���P���j�Y��YCF��i���Q� �f��2�f�u����"G��-�(���
}�@�=hā��R����bdBcq�M��S)z�:}ޓ<r�~0q�&k�eӘ�)bg���t%W��ƌ���s�����.!�g�[�p���_p<�o��}���8���@��6�-�L�Wf��b�
��Y�!ժ�C����W4�bÆ�� �Ɋ����n���!Q�δP<���0�5����6Uj����.�q w�:�פyM���YK��FO7�=������d�7��Y��4�x�Ro(�|"Ĩ�PY��@X��`U��)�w���$���@8(:j-7�T��o(��߈��i��A�B��:�/>�>�����i;t�S��A��1�ؖ��¹��0�O�
T*�p�e$��Y)7�ă'�������7YVve(���oP�&2��f>?�
x'7뢚d)~fٺ�6��Ӹ!ZgqK����NkTqDБf��p
�R8��f���;���V>�*_@st�{���5H���܎�md�]��{\�j��P���F�TPC{I�I���ź�J�ć�^c����f	�2]�/�]��i��{�D@挊�@��Jrk~���.�S�~���q�i3`ZX��*���hIH����K8�(�.��0ΪA�9C���ޤƠ��GT��O;G���1��݈Q�g�r��+�<���'�7��<�]Gg��Y3ۍ �PVS9}x��8�~��V�v��r���0w|M֠�뚆�꠯p�Q����'�4�mvԫu�NJ�5
iJ��Wp���$����)�~#Շ��}������5P 㪥�Օ�0&������c����c��%������וT�+u  �n%%!��۰/�u����V� �����?�²��呛9q^�z��Y��y��[��T�~���۲�b�Ǧ���Q�0�/`!V�/�d���G[}��-6��/!xs�jm�QX�f�~r��i�����z<��w�RcN�ί�;"�$x�=^�5ImZ�K*?0 �S�<S�:�'�40�7©�G���n\ɲ����
�:�l�5�u�H�wA�Lڐ��/�!w��C	���-b�G� AE��F�/��ݯ�6N�Z���<�o�l޼ՄܲCH�󙯧4a��Ju!D�&Z��yLw�K��QXh�J�����*�� `��\��4�3�/�&FO�	d�
3:vQF�M�%���Ȅ��^��'t�v�dK��n,П|�X�x�Ɣ�?�>B?�˨4��������'�/Z��MI��#�P;	�)\�Jj&�<*�mҶF"�j�k�ywZ�|�B��;�=�'92ibnL��<��#��j^ގ����C�%�i��������W_r��"Wd,��>��O���;̕�D�ۨ >���%O�#�,9ϸ��h`44�3�Cl�<��[p�����GR�	,���)����V-����G'	5U�v)*1���`�`�%1��p��:g��moAT
���bnw$��jؽ@��Iv<���Pf��h	�1�&V�?J��悖7������ �aP�S���Q��c��8K4�����!�x�nn.��(b1
��@�A<8��@� ' W���_\1f�O2��o�T����G@�H�#&߅�A��(qF��K�7:�����_�\kO���ޏL�7��Zh�ej�D(���W���Tz��]����n�	eG΢�pې���k&�A\g��"v�N��[��h�J�6m�ּ��8��b�qs5q�?��4��1�A��(��JG�����<�����8�E*��T��&�ɴkx�I�eP�˄y*Ǵcž�h�RQ�n�V�W{/�q��0�[��������/�V�`�]�bX�N���^�j��Z;��Ŀ�/R��п��mvv��1���=:���ֱ��Û�����o������6�Z���Z�l6[��
;�6$�g��}��A���[�S�)�i��}r�>�IW[Q��ϜZ��#=�]��.�0��`/���GA����8;[���p��@RBS�説���Ŕ�S��;I�C���#?�
��(��/R"�%ei<���>#�؈C8�rt��a)M��^)�5��5�g��ev^���D+��TOX����17�����q�zzi��٠�w�ѩ�U�=��g�%Q�w��^n-h�胜U���>/�����Kb4{B�7 E��E��µ����P~��X�����l̀rۋ٬ÈB�")�Z��޹]N��В-V[P�D��q�TT�q}B��w�g9���y��Lpd<�g���z���!���s�u�=���S�j�J��9;:�d��;C���j�XG-�~��_�5'����i�a���"�7��T���VU�l8ui՚�ۘE��%C��AZ �i=����W����\���ul*�#	�d�Et���@���b���#���4�]�\M|{dP���O97g٪�iFւ�W�=�8))�8���p�Y�~�uS�� Z���ǖ&�}
T��ލpE�<R[e8[�o����@� �*�_oa�U�@H�T0$\x��K�Y6�wP�%��N�j�>��JO���% �T�����Ң���R"�p�v�ܱhB}U��/z��_j�� �_ֹӌgw�;1딞=Nj/S!��T��qO����$��λP1�������>����`Xu�f:"]	�i��T�ԅ�o��7%_�����܆���4H�W���l��|��r��f߻�YoZv��^��C��SE���Ԧ�����p�����%�f舤���&4H��Q�*m����2P-����l�,����-R��0ei��� c��`v�]xԶ0ȅ�"�~^)5�Iz�iF)�M��ySY�f��w1�����n��"qgYq+>��m.�c����a��]�2��ntS&���8b�2$7���~�(�� /OP`5�����E�@���$z%+='P���'Ƽ \z�`y�TǗ1����uU�����(�߀��N(-9��Y�7T���T_� z:Rd�)V�����`�����'x�T� ¦�LZj���q����
+��oB���ɱ�:��i���7*��o҅��*�tIԭ� 3�^��*�3n�)�����m�l�m`�|�LbӼ��J,��,�*5X@
�Z�E�6���Y�b#��u�_*���="n�J�A���8�'J�Xb��s�Y�/��ٱt��h�S�ڴ��i���� 3�ٖ&2Wz��I�\k���T�e:� .^�n��r+L7Q���v���In��L��t:�b�ӏ�1ђeTc4�7�rZC��+5%w���\]��PꆹED�#h�^}�&<u����v
��,/��6p���7u��e��:�%�j�I���Kw�֝y:T:��C%����t[�, cya6w���>�����!n�]V		�R$.�[�����i� U�N9����0�����X�؍q��m�
���t!�C؎��ķvr�.��H��7%ӣ���-&�ν�ҹ�d�>0�W8�f��!Eo�1�iAHj�|�Q�D$�2|0�	� @w9_��Q�ǶTZ�������IS�l; ��C7�%5����(�t�"_�i�`��0��S�Q��lMcu� ��GR_���}e-�q�	�(ɠ���^���}�kq>���rv{����&���|�6�-�Ž��&�~������*�LΟ?A��ZݓT^Wl ��{�'�T����:���Q�O=}ԭ�-;�@�J'y
�*�=F�ݺr�"�h�|ե�Y�(p�1��jw�+��q߉���R�*�Įv�v}uT�L�l�깿I�"�}�U\X¨�i����%�c�Un3�@}�籐�`���m#�@�\��9����߻P
xF.�&`���L����:,���ŭ*ޣ�|y� ��T!c�D�ħ������$aX)Ȭ��r����c���߻��)��`@X��x�S��B�0M �b�[rL��Hh44�
"�y��kϡ�U��۰{)x�����U�RYTt��S�Z�b�W�x�\�W�q���3�J�gSL֕���}����(v�O�֍*�K�Abt?�-۫/lNH����S��J|�z��{Ik�f=X[��Hd}��qt�^�3�q����%ڜ�ZU�PJ�PY�s�F��CS;m��yv�P?|Ha����%��]L����392���u}x�5�L�3��&��hu�tA�,Je�d�j�L�ZC񖪌��؂m/�ۢ5�R=A9�)���	�e	��	 Z�s&@5�������)��N�xP�9�*;��2�Ѵ�υ�%�Q�Dv���Y�z��'�י\�(�Z���Xs�,��q��䴲L[D�<�@+�����
��h���@\�z��T�m�\[����$�Ф�!�P��|��cv��w?����5iex�t��a�,�X	��܄�cPS�J`�v?�f������VyD6���ߟ9FI���7Ξ@t)�@��4�V��M�̈́&P���N��J��م�^F��X��ο��M��/rɉ���m��_Vf	8r���({��%=�`�ɮ'm~S��6�A�9i�v�p
�����G>t�8��^�U�3�s�����1T}��1ڄ����|�Y��N&a�u��kNx�%�U�
�}U |9���V=���9��ҟB*��>�'�#�2�C˒���F���Gnٛa-�[���3X!��gf���]8�����W�p���{-n#����߫d�:��K)��[�2�\�nV-6��$��Q� �(�ʆ!�'BSfG��Υ0W�	��S�����āsД��<u`�WV�Q�����hG�ǰ����.y�J 6�]�*�"ހO1�%��r���q]�h�d��Mg�k����"d��p5�췬�T��u��慳��w�R�t�4[�G%|g䢾�������E�!��Lx���q����s/�i�aC�e����]D䣘��)u�����Ty)D�����,J�z���� R~9��n!�N�#��_��	����z�6�ЯQ�A�e�����Ao*���n�E��ŏ����!����-��G�]�L��,��9M��m�K\XI>a�t�[�k���w}JޱUy��eG���9�O��a�6�U̕��m2v뢢4"�]�(Zs�=�<�Mc�`��-K-D�/t��T*���y��u1��;ֲ
%�f�p$
3W�X�|�kgq�vg��QY���3�Ɓ���^��4�L��Kt���e� E8q�k����*�#�8��|Äζ��*�zt����}#�l����k�[o�qW C���ڈaW[���]{�[�K�%q����7b������@���
y���]��Zvsy/�UR�-�?l��(�!�4�S�O��͗���@&�
�`�%�t'�#����S����1ކ@vռv�z1���Ɠ/y�7�m��-b}��8����6֒ϔ�QɁ3��H�*�pFs��a+����:p?�b[9�h��[�}k{E��!� �A��ȩ�Zy\+�`j! A\�}/1�*<r�4�K�c
w<]b�����U-`�i�9�lP-i���%S4D�駉��r}�kz�{U��$���q����bw��� }}�1���5G�끁�h�˱LТ��:N颫kw��ze�aV��[y�c����&W�㈂�E��y�ܔ�M���Ғ���"_@Ӭ����Eh������[�hY����%���;M�?�h�OJ �	���
{��*�9euhO	N��^m�Ŵ�X9��p�
���O߆<01��v�G|ږ~M}��q�7����$4��Hv��¸�+F.8wzMכ�тB�ʻ>'�)YS� �-�s�4�f?�B/�5I9��A�b�t�-0�!^%� �;c�ڒ@24y҆1[!]]�X��f�d�A5�=ʀv��hv����Nˌ��W�<���6� u�66���y��?R*��"��Sˉ���*G`:����+�}�]|��0{/C|S�횫p���\56&����K��/�5|�m,f{���xx��E���PA�@�(��n!.K�W�{	@�|/ĢQ�����U�;n� �����,O�h1֛`���-�*�������LE��;�ٮWC��ou�pJ�D|!l8LZ��Lh"v�����'���V�F��S%���
�Ӵ���7�el���h�9�`�B��Ԇys�	�lB'}�����zg� �p��H�Ъ�z��Xy-\�+����fd�^���.,H�"��L�O9��N3�}8�0Ǯ+���Y���OaG��nFMF;*���"B"��AJDY&��':��##���Þ�i�C���T`>{���@��V���J�i���#�ԩ�g>]4��z�[�]8kǁ}>ȇ�x���`����zJc�;��DU`� ��CR��9yг�m[ʞ���?{�Z�j��?�t�ϐ,q��N � ��5KT��Q@Pk�!U�R�����@U ]CXbܬ��(�?Ƭ!
	��m@�<j��I�Q+�Q@Vn.�z��%{��Η����	��~�Mn�7b�3�Ք@�ܷA*�!	��#mu�h�Z� �
�5c�#¬���-٬�+�]܁��\뛻n�t@�O_$	Iy��lL���C���Z˓0mi>Q��Lڿ��àe�|Bm��u�[n(7��`S����|`�c�O�h�����e�>vj���GTe�!�Ȗ�n��Z�����DKe�^[�N�!��u� ʋ�$��j�c*9g4V��-��<�#����{��d8�vv9��q�y��˵uWb�4$Ź[7N
��Ap��Z:22���m ':�g�����S6R_'�L�����ȟ�1��������y<AD�������iD*�0��$a��ep���5�ДQ?"�e�G�]��/��x�혎v��q��)�
�S?��>u����d`]F����qs�h��}�r/�^��Mw5"vzi�{���"Zǉ��U9����Cl�X2�D/d��ᴟ�z���َ&�V�]5�G^cZ]tR���$�ĉ�dO��YD���<�>�X`�)Cʧ�����P}hsܔ%˿�@;���TZ�S(�5.1�c��f���g ��]����$����c�q����A����n��$�=���2tu�+��4ƻ=_��j�w��FN���<�*�W�94�G���ieuw��OP�\9tQcޒk7C�1�6�h�2��P�<}�Y�C�k'�s1��s�0jϜ�ؕ�d������Y��) 	0yz��tJ�m�0w�����ġ��W����`�Z�۰l�t�Pn6xP�@p籗Lf�l*L(���D�3Еe N�_!�/��t�x��&I�(�^��IS���oT	5r�>��H ����F[��z'|f��̂��S����[=�ڸ,n�H �����f�ܷMz����uagG�3vs���k)ř;��[W������ 	3NT��K|�M9Q��j��X�آωv	4V�v^s���M���ס@�&�ѓdDT�U-q�����Z$ds
��_��o���ѤX0JqO8E�����\�vM	����h�î�A�����{�3�;��)��e�O
�Mu+E ѵL42ޮ-e���(̼N�L���J>�G���ԭ�aL�1�Hlˊ�~iX�K0�SR&�=�s�g�&;SڣJ9M�*�d�O��*XM?����E(�ÅS*�����b�B�%ḱɌ�s^Y�JS������}�P]�>alY5�M��x��z\��O9��oeD!w
�E��?_�&,������R�i;^ݣ�A��o(CȈ��=�S�D���:��F�u����y�/O:���|"��hsķ��jŅH�ŗ>���3�YA���3��A�$�O7�"Ze�٪�BM�A�[Z�p�p1��Lz�w�t�Ek�7��1���ǺP�G�XĶ��*c��|�u��_ɂ�d}l�R#�h�����,��-Ƅ�h��;��{b��|iS!z_����6�rg�L^Ϊ
�ҧ����N^TK;V��3�[g�O1��*����!J����(����^@B�2�6�1?A�9s%��}��ċ?;��ƺ��ؾ�J�<��q�۩M���F;Ѥ�,�} 1M�@��h��+�h	���t{�����+���#p�)c�H�KoV0#�%R0ѿ2��Q_$V����<> 9����>}�w���ko<lΦR�x�"�{�k	o邒�\}*_����$��)!���2�������ɨ�Uc`��G�{>���T��|Qo4/}�zH)���ˑ�:�k��7L1��WA�A�!&.֎g�D�է����PjD��ޘ$����V<Ye�Y��M�S�r3�B*KF�0����6�Q������K��8��ߟ�q��33t3�C��@�ٕ䩠#�U;�.R��g<��C8(l≾�D��V���K��;���i|+7��L�|���.IN�"��]�c�N[�O].˿��o��8K�ĦD�pA�)+x �A��%��02]���V���D��x$��SJ����K.!>���o)\V/|.�>��g(́li��~h�\�6��s�G���eڐ ��M$��P��*��RBO�\�����٬���N8���$�3�l��g�q:�����J�~t6^ﻗq���~'n܎��E�@�sc$��t7���)�h���<�a~���WN���(o93��(��z��XL4�k����U#0��o2�!8£7��.D
��n���a���zT��*/�X�B
1&puᏱ�D�<77�,\����%����Ů��Y	�Ђ>I2����ɉqޟ�L���+V2�h*"������o���Ɵfʆt?o��Q�H%��]%R�-B~x�ze;!�n�{���PR�q��vO#NWR��<D��ol�e�WŨ1�	�`�������@�������[$�O�v>R�P���¾�C���:m�cr������E�~[��J]T�>ү�r+����V�5��_7�:��:s�妚�Jt[*�M�o�yˎ�7�0�uR�S�]ıRpQ���`���.�&��5�	�M'$�_"�p�r4lv(��"6̧}��Ggn�U��O�Rp�� <�t�b��(Z�^�Ѷ�\VVY��'��}֣c�����Ou�1����yO�BN�ƥ*�@���XjjX����4�x9���ėSb�a�j��k۳&#AR��A],6p��{^8��d���iיV���?91 ��U'Ί�� =yl@D�߃^gQ�'��Gu��Z���o�W^�}wZ^0D��,	��"&eO�LY�ܮg&��+e�M5#�#oL�$������:\�+�Z���q�?R���i|�59\���d����d$D�ޛ��4]���(#rn�$���t�w�Y���$�I����R�a���ۺ5��$t�ŵ��wO�y�����������5�<jPxa�dn���;2�/���ɛn&#���f_Nך?�X�G�吽�z)���a.�uڪ��[Z�Y�\{��פc�AţJr�vBJ-��O�8V�Է'b�r�4饷�CgΣ�}s<f�Oo h��7_;��x�c鑧-�u�1MrIY��RuҔ��x����7+�� �Ne.�Z�����7�/�%�K��%�&�Q��7J��I��s&�O�y�(٬[(�}�ݾ9>.8����ٸR�%ݝ�R��c�O�X�3�W�|�O0��@ߢW��X�������SР<c{J��	p���@Iw�j������clfo�[؁�n��������Ws�H� 9��{�$�eRA����~��h�
%��*�ʍc�Mi�5ds����c��L�Ku���	��:/m��k"�P"�@��	�Y|l=s�RF)���Շb�s��~���� �6��@[��Ҍ�%^�� ������M%�@��j(�E��f((�����6]��M �����a/9�¬�g�Un���q�^PK����J�1ʞ�<u��h�Ք�T�@�Ѣ�uJ�h �c�򓪟ň����5.�������y�%�X����d%	v !�4�;��d#�jt�j�4���^�E�����%)
v�4Ȑ�2��ҵ㗨q��F�ؕ�T�:#�~R���햔4b��bbȿ�Ek��Z��aЙ��0ι>x+�R-��_��l���#?�$�i�h�N�:;���|?�1��!@]a������\%M��4,v����χ\�;�4aqkS,���)����$��n@�N�7s�MY��n42�W%ȿܒ�$C��	��nAC�bM��h��pm���õ��S(}u</���/h�=�4Wc���?�XKk�
��n���K��W�841����g��g�@0��[�m�1�%�-�0SyN gB�H�,'�y���Y[�bg�-x:��B���Y��Ia���)���gr#O���__��t#ұ�5"�J�K	)�1�T59�TiI� ��?J�����ɐ��(a(=��;�O�8�kА4��¥�ա�� ��_�e�'`�Q�饤�t���~�[���!��/�'��	'�V]��>�\�%"<��}''>DG�<A�\�H������7�\6l�O���;��.��c�� y�����~��0�!�m �����x��,�CS�Ůs!�Ll��缆�c<��ǖ�5��Իοh[��'
6;�P�4!&=�m���R貪�h�n]w�'63���EQ����r]R�M娎)7K	 v���%5]/O��{`�����I��D@+��xM�����#�	U�z����&���):�㤇��A�����
�(\��:�"�
�1j�[�n�<g���iE\��ۼw�9�������0Y����;�V}���eZ;<{���\@���A��p�@{i���MS�>'���L'3������G��Q���+{�o ��0|j�`4ST~�������׺,���K�"���*JpéR�Eϓտ�����������1�&yh���fT�FC�xCC�ݲ�nR�R��"S��P����7����r��QM YP�a�nx��3��m�=:�?�OԨ
}�0#(��O픋��um+}�lRGm�e�sdZ�h��)TǭI �Vo�G�5�+�b�t��!�	 ߉zI�p�'�*�g���ʋ�֎~��{��hm�-�U����S2'w�����1 �����1aA��+���ʶq��x�U^b�����|l�����f:b�&Z*�QVe:�W�9����pڥrO{!�BE����6wҁ삸��eҸX��^?���ͅ�D��Q���~,^eg{�����Z;Ũ#�w�9���i���UI�oO���;��K��N	�$Zb���?�����]��]W��B'7��+���V���v���ٲ�j��2))iy2�pީ �+�����"!W�ƕ{>"�e95CBz��O������c����<ְe�F���N��x����U&��7�Yz5�&[w��S�͂�~�z=���'�$ZZaDG�6�~w�)j���T�a��RJ���Q�#����+V��C2�)P,Q?��$A�Jbe.�yo몑8��Fs����[g�Hy�n�y �����g�g�[!�ee��F����y����毷G�!9P7��e��q?�=<���}#l
)�ؾ��%���#;��*�mc��њ�&���j���1�gD��eVi��4w� �)d7G�c^�J�]
������2>1�L^�7L#�Y���&�πh�}%̵=o�Ѝ�/}�uZ�"><2�h��a�D2ײn�Z_{/���>H�K{��,��"�"�Zs��]�ױ��S�r��P���p�tZ��������N��<X��?[�jr��n�8�0W� h�O\��aΡ�f)Ř�����!l�"����1-�us�$��?&������Cā.���32l<�����I��x��׉��v��XU�Q�:&s/NM����9"C&��|;��Q
�WZ]+/�gV{�uJ+�Vv�F�Md�;�0���N��#�L4� Ti�������Fe���w�������'�F�hk���̣<*��X��?� ���2*�}b���>;F�#SM�T�RX��n;�{����>�6/T��)����sZBu��CANlc��� �U���!�|�fEt-�Hd0�'@ Q��X] �=g3}4O�m��w�� R[�xu��!�zZ���	�h���#��u�gz��=�T�/p�D�����Jo���=%\����zUC��n��΋��U
$00�˻Dp|�����s��v�kj�FN��?��FtV&�4��KgR���~�8���F�ۄ����zZ2Q�A�ܙR#z`!�'�ԉ�g��{&"�c�w!]V?�_$�'U5���H|?U�}]�#t��`��Y��W�Y��M5sQ���4i"��BM��C���f.oc�-d1z�ZTF��W �	2w���b0�����`�:���S4̖��U�H�����~ѐ�c�k����h�n�'I�yh����D:d�g�:-ʡƇ�621���	�\�m���\:��8C���������*XRyZ슺^	�v�B�RU-��¢��&b�H�g۩"���s�֜�v�T1�w�b�!��(��n_�.����D"oJ��
+������}:	�]6�H͠�+�q��(����^���΁���n�w|��<Z�<��E�|��laE��$����F��w�|���o�Ԕ��"J�h�ʬɑ3�1 ��ĸ���naY$q�ϴ�#�F.��RS���a�_Ye-�t�C.��(��_��6�[�u�A���y��3ֺq��AqC{E, :Q��F�6��w�]7M��|?�!Fz�5��}��n�A_�נ��ֶ�9+e��X��^�;�	ݸ�
0�?hW�*�
²�j
�C�/����:N�~,K���o8��M�X�r
�0�CDF��:$1I �����:����ĵE�(1O	ӗ�K�JB�w������.c��M����J0���JR���_�~=`h��e�Q��?hjjǙY�L����H�k��P [ѽ� 1�G/�iN�G��ݘ%�	<6D��g�9�v�gr������MZ��O�N\�G�Q�����۫�,��tz�%[����t��u������6X�a��� o�$�L��Tv'&�����(�*�n��.x�)%0���.���\�g��?����o|���r���/AR��64��jLU��ӿx��"8 �4��wG$5�"�BxOB�5��������$S7�)Զl����U��M��¿�����?W���Ջ��|��ͥ��t\���kA�$ܧQ�`2����]w=ݾ�'������??�ՁAo]jGgQ]�7s�tAˎ�ȭ.V�&�:�M� f`-;p^����z�5V�=�^���%D��
,����'竡�g����4��饙��/�4p�%U#õ<ov����^��O��pQ��FPD������'�cD�w藣j���X��z�.�Ygsq) ?s�-= #;*WF�����Kd���L�-Zٻ�Ѱ+` ��0��� ����E��c���Af��� ����z��?����ٯ��\x5���ߔ������f���|'��y����`���qm�Z��?�t����yf�Ҁ�X��sZ�G@�ս<p���[��?s���F�W�L-Ca���?0ދeg�~��P���|9�X!}dP=�M�2��,�Gq ��ݡбZX��[����@�LI7E�N [�!��pD��x��s,�\�&�C��u�ڗ��Mfޛo��H�����	s[��O2��gww�sl��V�	�~t�m�zg�U�ӢU�d ����[�y�m-[��2�}qX�U%�v雫���X8� �2�q��1�r��m�0�CQ�R,���.�#l㗎Z�ɯ $~�Zj�B�F1EG�f&���5އ�@/�=9+jf�ıH��oO�=���~��"��qq�j����m�.�>�@��O��i2_��w�j�h���3���{�O:��ˁ���H�G�z�Q�k��*,Jdk��1�-
7�S� �$rA�UG|�4Ď��'���?�t���i��Ik��&&�O�����<��;�*���Ap.Rd>k�+C~�`Ԑ<��EH������.d���,N��-3#\L�

��I.G��
]�ϰ��Ak��,�D1�ܼ�PSNh@����i������_�;#���W`.��=���<��"Q��$��OAN8���x��������c�.$��ch��[q����g�v��?+�Q��6Hc�b����7o����9�W��\9rb���{��+�U=��M��r��]���H��;ɶ*C��*'�\?L�U���Bhi�q�-sr���3��Wx�;�B�[o0Zʰ~	X-�i��ni'	|91���f���)���7���[�ч_e��.9��y,�(�E�y�ܸ?�W�	ԛ�v_�����P�KV}NHHۭV-�ĥ�9F�T� ��Ɗ*,���&�7�G|��H��q�dbFM�T@��7�(؁_�D,��Vd(�ڮֻmÌ�*P����������W�B����6g���鉙;�l���Z;������N�0:U��K��":iI#-" 2��?��͉��س��D�tF<��/�nӄ�93'e����k�;�e�h7ڷB�=�r�n�HK|l0�~ �1� ��>�Ί׿���5r�m��5����A�$&�^
�Ty���M*~��5�~y�����8a��΋�;�i�2P����,�.������%��kI��3/L�����"����H�K�:���W����w��;-�d����Hg�0��M��g}u?��D�)�b.����J�������Σ�#|�� �*�"1Z��O�����r��_�g b�I���/�nC�裮�v(0�� ��/����%26yl@y_b���pY�cZ�Y���WwS�e���	g�2��v�]X8�	M�ג�2V񆌚[��vno܃8x6GTNk ��+��K���Eñ!uq0�:j��}���!`X���P��|�u��zF]F:�,���SE"'���:����XƟ�,�ȴ�`�aD2$H�_ɟ��m�><����:�s�o~qK�nsUmd;fd��Ѯ�$��.*�Q�Ǧ��O��I�y��eoܡ�F�d�lr�m򣲢DR�B�����j��I�@/9�,�A�|��\5 �1{`<1	=��ǔ��H4,��t�t�Ǟ��c�g&���E��>�9�Ɗ#��Pz0~��˜��*�ģ�[�7C���x�L#O-�R~N���t�ӏ�*q�o�LtK�Yg��)Ue�#�X��k$�����/.��w]x�8���nt�.P^�䖄k�_�i_��b�+i�@\��q`�S�ş��ͫ�ԎA���_��Ϫ�� b�O�[6H�=�^\��j�R;c�;�wH�\�XҎ��}�C0.�)���!hKn/4�!�'O)6���MH�<�,H
t6�����V���$e�8+84b�U�.�}Taԥ
�f��^EL�3�!{�u�r���r��36ji���r�u��1��s�#|0���ʅx��[߄���	|e��	j���SU��}�AH�#nu��)]y���n��ZXE�m��$n̻<0��q��f�}I���PӞغv��Ed�͢]�?@XX�ʃ���ψn8^�o�OR+��*��i�<�V*ī��i��+EO��������Z��RD��ɦ�*���D! ��JN���}(+a�����4c�}T��������,t��fK�2�g���x�BVƕ�)���y�}خFO��M������d�kD�b��F��8�v � M�D9���q����4Z�X�0a�����Y�� ��J�����2�s�%̵����wH�o��0�F=�+�j�u�����!��)"��l�/Q�$��C�{t@�m�7�����S�����w-W�*�O
*�n�3ok�A`����)j-W���aK�CM��u~���y)�d0�����VnT}ٌ'�W�9�� Zc��=����K���kr�T���e�y�����̣�F%w�\�h�瘣H�`�ͽ�6�Ql��F9�̬G�z\��U7� �r��Pkד�=��4����5='ӠJ]A��ߵ
��k~m@UгZx��ޢ`iIMP4�#�V���R���C)pwC�8����@x�sNx]��M�ՋԜ���Mb�g�������7�^�zۼ�^yj>�ΜɆ��R��J�Rn�m�k$&g3�o���#3��X^q�����2���א�*R�@���*I�
oG�j\ཛ�ݾ�y\��Բ��Az�1���[3��))>�=�*���axr��סjA�x�o�hf���?h9�����5^�"���D�q�� Wѻy[�N#s@�N�1d���QG���jpm ����ynW��ߙ�cq:�L�Y�����!u�or7�*n�^5\����Ka(BIl1BW�8���]�tn1�2M��OM��"M���E�g��%G���s:�����ϿS6�mH]�Qr�H+Z�M���q7AЗ�����ox���BD�M<����gE��3��eևC'B�v���7�F�ߊ^{�)�`�P
#�B���
�&��u�7��g Gl��i3���˷E4�Q&{�Ӟw�^��Qvm1�����Ǔ[5wS��e	%�K�w�iR��Y��S�b�t�/s0<CR���!+®.�'���lq�Q2N|Sh9l�>��Xc@�dd���'�iF�Cl>�C��K���$�lƗ3�htȝѽ2r^3��ʁda�����@�-�;%����mk�=3:g��^�����̀�u0�5�su�������}WPI��`{m�Y�����^���z����GlM2�F2�(Yj���]�m�9�R�X�0�@�ypr~���1C�bkd���,Ӄ6����5�O��T� Lud��~n��y��@&�H�%��`:���^��7����#V�.Ӷ}FD:�A��l[��K���D��܃)��;|I*-Iҧ0
R��Af\���d��/���p�s���x$m�);�B>�n�e��Ȧ�_�	\Uȴ���#=y�;l¨ ��Է���T�t�8�9s��,��N���B2?�/�۱2��w]Y�p��|;Y�A�W�!&����"�MS���?^\�d�[��G��H�jB��{X��j�^da��D{!�4b����8�~���Ǹ4t��J�E�K�f����[�'}M�з(ݴY:�Z݋hj^V�%N�a���S�@������_#���cHI:s3��O[�u���D�_�|�L�(��,D�xm�����I�m����@��L;�V�9 @+YB�h��{�R�r��d�A(��0"ٺ��;�(�z��{���=y��2��՘��@9�M���P懮-�{�L�jkAI�#.�a�l��h0@Q��,FB��X4.�^8�{�"�hA)Jh�%����XS�:Sφ�Qth�j�������Q{�em�=Ye�̞5X��y~���V�Ɵ�}I�*����uYg�ľT�4��m�� ��H^s��8CC6�':��%0U��ۥ�ߤXbdL�mI�]�(��]�od����[LWs�$tgӃ�ἋSL��������p0�H6��sS׻]y�K D�v��S���f��k�m����ϴa���ZY�!�n�����p�M�e��N��4��q�y#8�5�n����PӭlD�B&p;h�]"�U:C�!p�!�%z��U�Z��R��Od�ދJ��K�o��c [��F��k������i�\��B�Kc)�:@[�W�ZH5�~t�����AW�����������(��ACy��{a�>��q;�{e�%����J�<�/ �e�L(�������PJ�����p�U�O�{�$�Dp��x%ij9�%P��=m���$��&�J���q�g+A�#4XJF2́�*�ձ��_�z]��p^q��k�m��-���27��6.G+���K.�x~����u�����Ԓ1�n���]� _H�aǝGG�~������٤D�%w�N���^|�:�ځv�G��38�1$�t�3���o]�#q��C�N�;�zWW��0E���>� VK�6O慛�R~�j�ɏ��I-�ۑ%��I�k+�v#^sֈ��H��e���\=#Fb�D��v�����!,�p.��޾0`&�'��e-�y��Wo�Rm�K�Ę���"���!���.�=I@�X���"��H�A}-�?�MBᱥ�������:�Dp���^99��t���1�
���5�Mw�@��p��W�z���Krlg(ɕAi7�0
OR������:�V��vOw��m��x>8�Mi#��v�Mh����I�k�Q���!$`]!�$k��`�3Fg�v�& ���H��G,��~r1��'���r���D��OjĊ�����:�xb��.:(o��v�G��[T$SW���:��K���/v�+#�W.qRk/٘\G�CPsFݼRy֔|M��D2t�m�F� eO9&:m�N�����7rs ��CaF栐���%���7V�;�φ�f�n�$�x��!�hC�v���8.�%X�\�gUqa� ܐ�-����"0"�찄��.*����"��3���W�%�r _)i��]O*�Z�A_�]�c!�p�+�D��=�᪯��9ՕFho�?���ط��em�����q���#�9���:O���Io�����i��[��}t�P��~��U�N��� g�ũf�1�Ӫ�c��>�L�A�o�A���Pw#�M�qd�h.���v=
��6[A���[�n/:�q�������z�I<ߖZ�ߦ��_��ȼL=�)���Gۉ^��u�Hu2�O؄7�V�|R��S�N|8��,7ka���D�ϏPg��� ���%.����%dJo���(�����T���D���\ք�W��S�k�;�0�j0Ҩ�A�]A�&�LWU<�y�:��֞ ��g�o�F �"�F/�nNmxĊR� یկ�Bt|A+�;��&�nŪ�mq�Ȅ�����\a�l|`�`I��D~�����w|��n����6�z��8#��oR�Nu@!�UA���Hf�su&�O~lN!iOar��L,2��������_F��^���A�^x��F~H�eɉ�*�}K�-��yA?����^
�7<��*h�ꦉ�5����i]q���O�\�!&�-��0_%���F���Y�a�a�S�>J9�oh�/���!>9Y�F}3D*��ɱ��:�YTOoۏ�;��`�����-���7��#\=1���|J;��_��^��뎧|*�Zo�RwM@��(\nNx��o�Jܴz�k}�%��ťsa H��J�C��4�ԿM쓌�mKz�\y�p�8��mGR���Y���4�6��+�1��z	I�3>�m�`n+|kN�qUv�Oרa:0?����AD��޲e
����3MU��e|��ʟ��b@˒C5 �J�+pm�
�z7R��0e�-��F	����7���@��
n�K1\uچ��lD�EM��;x;������|��æ1�V��2	�Cmc�|[��X�[�� ��[���4��:�'T��G�_Q�)���n�o#�֧7��'�GEO�]��D�;Aq^��$�l� �̳�����^�6&并�{WdUyh�qAS崤�%t��w����~�fq,���8�� ΄�S_��,�?/��E��W�ZĀ��wN���W�Ez�
�x'X�/�:�����A-ǹ��q+��Ē[L�Zrw73 ��ۏ���!}��=�ߔuNٯ%k%tj�|AKe���5�G�뤹��B|Ȁ�>���q����6��+���e�n��࿕����Z;$}�%�����j�6���H�dB���pO%*��'9O�:�;�93�Qq��r«唠w]�c�a�T�"ۜ~6��B�C�A�F�����î
����:>���s�\2Ɓ*��[Q4R�OV�@PU�V?�/��h��vj���i$Sr�\�"�k'vbk�a���s=���	��;n����P����
��ܜe���fV�%s)�ruٖ%-�[Z˯{i�1�T�#=�u�4�{S)��y����=
>��I���9�z�[PҌx��C�B�5��@J.��M5�d����ۣ��=А�[�S���'~H9I�/�;a���>W�6�5��`���Gl/�o��ѧ�=?嘔�]�% ��n�U�0�>Ǵ��A�n������!Ror���^���}p{t+�ȕ ���}�oo��s�RK7�a��ٵ>���|��M�y���U�6"�&��+�Y��q�'c����X�-�݃]u���tʧ¶���FNb[���*])�]�����c��L0�᩽D�u���/@B5s��D	�CK�&�W���*��V�`r'z�~�����䆊���AN�w�l����Hg�i�x��<"zC�h�Ŭ?iB�+}�G����;Us�`>�C��r��� Ŝ'= P���4'
����n��Z,]���O�ѧd�O�C�?����{��Fa����(ƶ��uY����j��E�������~BV¶mJ2���mNCAYK�@�����LϏ@��i�Bz��edY�t�e_W�m!0�=*J�J9u}�n�x��¾qg��?��<Trp:�~�K�`%6��>d���+��{F�zߨ"�E�|Nu�~���u#|�N�S��É����K��#JU��
裈�.���
6�v�4�m��IJ�m�_�Hh��*�������7߆*y)��4�:����۲�S6͵�>/�ǀ�A�r~{�ߟ4��p�LY��-b�9�.o2�>YGDTk��P��@'���['U�Qޭ����}s���t#�n�w�r�r�B�H�" \�kC�Co�ޕ'R�@��dy"��W����A�B�x�b�U�R�j���~[�����Wg���-W	Y�`\����F�e�h\�0+�84;۸3t�7���z��&�d�u�h�dT�l~���z����W��$�
#WV|W�(�@o���3�H��>��z�;¾���	�A�x���Ss��[ َ��4����s��u{?�SD"^)*�DEb�H\X�|y�Y�!`5>_�������Pzu=Hޖ�YB�0��8Ѥc� s] �߼��3�33����=���I�tѣ�#HDb��r�y�,N�Em��X}d<a��1�0���@�-/2firDp���}�֫��Ɓ�X�ڙ��-1bI��E��/�
��^~ys��x�o��e�����g���_}�x{�\�֛��f(]��rt�4�Avj���ll$�q��͙4����d�q@�����Yf)ny&W��������|�A�U��s��d�x��5E����c��N�g'�4�۩����pb����Z���A���b�t�RAч�m�
�av���X�
-��86� Q�gFb����YՂ aΧ��O��Q�t�]x��(L�������0v�>8lն���z� ��KX�Vy11G�<���	}hz'�;�������x	�	��Z�IJ�0�|���o�P�G�AU���&!�]8�8��%�V3zW�{��(����7V��%�߁S���͇O�ne��4�a>OB>��KD��G���b���� �'�x�N�[z��j�Q�܄�6���6,��2��g�i�]�aQ���uX� l�6��"w�8���,�a�#DUԌQ�Pu�C�b�P,���[�ETt������t�����]�uH䨛8�9 ������/�q��?�$
��2�s��R��m\ea[�\��2�\��6]QE�ߝء1+\�p�:�oZ+DQqK��i�����au4^ݷ�|sYJ�V��������hO����4-f[��y}����f$��fJ����b�x�c���87(X�]�*ԬƷ���J�U��{F��O��,�iy���ε�������倯��w�� ,�sf������:�rs�Y[T*o���O�?��=��÷~��o}Xb�MUp&��O��1��EĹh�X��C�sẞ�;�"Z�[Ns�k�Y��Z�B�(R-��7
{y�tڧ6�6o�Epk���C�?�b�| �]�BH�\^kv9$%Ӱr��������w��æ���N�r~����h���~b�w���tU_DC]���H�+,>�I�ɀP��>��l���|�u�G^r�t)�{�U�|7�A��K��������-���ɼZ�'N�nҶ�c��~�j����h�{��yb��f��Y_8;,�y�C�����o-!�n�MՃ�*�6L9���f����&�_���X
I���� ���ɰ>ǗRq�};�j�)q������J�OW_�>���8�QMFt�\�5�_���0����|&L��*r�DL��»mS�R1����YM9�y<g��`�.�j�����e#J>��i�׬��J~���II� Ά��-9��o��
�����W�༭�I��m�}����u���!C[��S?��@��;��v4[��B�^M�^���+�i=�O2W�b��\������߮N��
�m֌P�o�����!(�}g5���kƹ�:��}h*;��R��I��z��Z��-[F�[ǲh�R{�+��X>�xr��R̴�ɞ����Ã����4� D �����4�1��%��V�-��s��"�oݔ�lFU_��o�5���f~��N����g��Yl��m����f3�Ͻn����yRm�6�Zc�����;��������*�"h��)��JxŸC��ɗ8��P)�}��K@p�"-Ve'5'�l�P��C ��`n���"/;
Ytٔ��R���1������Q4����y�̥nh�IA�� ����l�C�_��E�e���(A�2%�:���:�_���NڠI�O1��H� �����Y�թEU���[k��7��g�.���:M���q`� u�������99o���fd5���i�x������� �D��[�N�V�CTd�)�v����W(F�-�<�zaE��Y��\��냟�ˁ��^�~��O8�I�dg���l�yhU��^����q�{	��q�@���濛p�xsf,AC�J9Tr���O2�Pڶ��d¯~q��M�2�3V荪b�m�GCQ����D��mB,�U���x���r����{�#��#7�:�
WI�ԣ�xS��β*o`��T��D6�
�"���?����6,��r$b����IqT<+&��1��zr>�b5��a���%����0qI��~�hc��R@,b�	͑�ָw@:0Bt3v�U��@"�Aț*�[���L*� �lLB���hc,�DI�j��B)>��#���T�ƫ�g��}����=�ǀ+=�#�/׈�-�2)����.�]�K|*�.��_�m_�Iq#��i�B-x䄂5b$�x�:]�FEY����
�/sa�^<�Gv� e�|�����6�k��m��^|�:R�v��;�!nN��j����S[k�o���y���/c7�dM~�Iڕ��sL�����\��XQf_Ev�A3�n�ݫー�:ӯBp!�6��Y�.@S�v����~�,�Y'!�����@Tpzgɡ���I|xg?v�׫\�Z���9��/���^@SHb�]TT�4O�g]ܞ�;��Dx�zO=�$���,��ΰ�
��Jܦ�)�T�E��R]W9�Ed4���&dC�)�
�L�kl��3��v��t���L��C1h����}������+�,�4:�pL�[a�$���I��a� 4�-����c�z^^ʠ1=���֞�a8Ɇ�#T�;�G��!j�`_��T�kIQ��ša.qI/%��ŕ�$�cVϮ|\����]��k��O�4G��F�~�s	S  ����Ή�U��6Li�U���<ēqTY���UǛs
.$���`��h���8*���	iF�G��2�NvF3�=��~��EP�-,%�T��x<j���{�M���hw��7��?����?���ަ��@GHp����ng��s=�6IG<z{M ���� ,���~�	8�)K��7y���GFҩ"T��T��7�ی� 7P�sq�C��c��\1x%��fymC�� �=���
��T5xi��'��K��6��S1y�\'�"�=��~�Fh�������k�9���5�w&YH�b�B�!�)� #�EX�Y�Y`���9�R�d\8�y����P�^��q��l*��4�4�?�^$¼?^2�#����F�@�uH���O�rj�]MW�;�)�*���}dyZ�v,�=������N;���_�0}<��*��������ᢅ{�1Iy����{��!L k�e�m�[6�?cv��n�<L�����Xr���y����������Lɟ��q�	E�`
��crUP�$��A���O���bS���M>c�X~V�yw1�����j ��{��(��&��S�c�_>*w�^ C	WF�|=�E�6bĭ{v��`>��؏����*�����~vȺ��G��ʗFB��q��a܃��ּ1K��lX�p��3ZEVS��!�j�\�J����e��3"��٪r�13)HZ��jN�}����H
u�@���"6���{���G������x
֪�Ɉx(��u� �|�M����@)4j"ఠ��?�W|��
�9�x*��"�8F/҆Jw���c�k�Gh�)��s�'���[�H�����آn��c�a(w�[���4�0+op0`C�h�)��d���f��b������:�gRSX��IWT�U��X�I<|
���lJxN��ilIԓ+�/P\�J����+c}S�c��
E`q}�y���`Q�"�N]��|K����Gy��d����w��w^]z�<\F�Ι'ʹ9�쎧���>�,\l=�'�sT�ه��x��FWÉ�3/n�5�T +6�������[.^&���]����yA)��C���s8�E�7%s[�xO�n&�[����4f=���7g�U-�X��P}�D�>G��v��)gs��l/LM�U��gxh��TU&K~c43^<5s$�϶���ܩ�����.)���=z׈O�J�6�O[�ww?�!��(�~6��Ă��|KuG
�k㝡��+����>�.7\m��*��eM�ص�_
c�����S�v����_�'D؝��q�D�<��-rvXK�TX��pu]�2\TgD���������a����*8x�S'�(����/��3��$���bZۂtM�u�ͤ�얔�q9os�-2��2�yŨj�� HH��н�,��y�8^U�P����'�}��3wl�Y���Ik�<����h�?��l
Ē���Q�X���p�@�t\����1�����"�����2	�������7J��F��5K֕��LR������[�����2K��sz�gn�!�I#�蔃�6Y�_�L�ׇ*�59`�y4��M�����B�j	�����9�
�һ��wL#��>őD���͒:�\�xN�r���r�F��<��c	��w��c%�%J�l*@���ql-���"�ϗ��y�F:�;�C����w�TBu���ͬ�Y�<(�nK�K5��Z����j������n/�k�ہ<�{C:��)t�ߐÕ�0i�|UN�^%��_� ۳���>S�)�%D�*h����p<�w���Ŝhl��:Uҩ����K>��K9�{�W��:s���#��pH����@��T���/����C���&d�!��5m�؝��<��uS�p���p-���ͅj�C�Ȏ��;������
N��[|S��V� ��8ƿ�-g �[�N6���2��9�:�a``��f��k�e�|�K���$c��<<)�k2~^��IZQ#	3���T�U>�g5P ��c��q���|25���g#ϲh��zOb�V�����e��rɿ&�WB�y�)�ˈ���А��$�B�5*/��E�Zْ���έ��p�w��8�)O�6cG��Zr���j/"�g����3lith���ζ,O�&���Hۀawީ���t�_ʹ	�<�$�����ه+r���������_� ���h���6���.���9��i�ax���z�ҚoR�A���q�b=�}� ��.��S�Ne��X,�&�
l�
�s�7I�6��e��A_s|ΥJrZӦo��C�(���e�x�r��j�!�rX�jq�&D�=�s����ȈJ�C"P1+1īlx)z��į�C^���=���ܣ[�_���t��������戀&8���Y�!Z�0ܤ� ��x�T��N�|�"�G��<��/4�ɔ�$��v��JO���k=�k����DT��C�X��tW��'|D:�����3B�J�!�i�s7g�GnH̴�{~���^�oSݜ��$ξ�t�*�-�P�Q�@<Kӝ{����7b_@�ɍ�t@iw)�y�<����AMd�Zo͈���S\d��ho��#+Կ�9I^���n˪�a��̲+7����,����6��h�{�e�/��=�lo;~nY.CwL���*�O�㰴�+굃�`;�a��5;h��e>�Ng�	(�s�E�wb'U��0	�{�Y�Ơ;�5��/�(r{���L��=Q��u-�yZ/o��L8Մ�R�c4���s0�E�Qo��J��E��j��`Y�%����(2[�c�;�!@����kN�bf�2�����ƲHZ�ߌqRU0���ջ��Q�"���l�^�eF/m�
�TK��Ӯ���AN�(�-��Z����ҳ	V��k�}f�����l�3��S�A��M�3��Dj��sd�|~�%p�F�2AVE)�e
���z!�wL�ꟼ�Н�u����Z"x
��u��%K��rh�������j���T�� �;�{KQ~"!��F3�3�RN�Fy�����D�Fw��;6��&�ֵ0��8�<g��T�_��[� e��@�F��C���T��~S��$���We��$���cSn�n�ǝlc�a�䪦�T��Lh��X��b�r̼X]�{q]�4j-��&��>��8Шz�`�i�ΐ~[(��I�w��po�y���s�R1+(�+���,Rc����*�<Γܵ��T�a%���@$��<�b6��f�䩕 ��ggp�geRe�K'K�=�K�r��{{>Ŀ��>	�憦��i�����S���h�
���v&�7z���n�5�MI�g�֒��-a>���g8I�_�p�n��]����g[�B���O*ګˮ�=�����ؐ���0��{рZgo��0�ܮ��v|4
�
F�2P�Y�Ԛ�r*�g�<�'��M=���bx6&�X�S�7w�>��&+(g�J_&��O[�x��^V�J���{;��i��V	*q�����i3WZȗ��2�$�$���F�ރky'������� KUs���!���2�q�C�P��$.&�n@"&D���!��g���B堡����7�xa��U�K@���2)�?PDG�� u=�<&N��v��,�>m��[&�wc� 0�-#a-��,sṠ�xO<��a��3UW;Y���Y�fps���n�Oz�s���gqzD���F!���I�]�3[��\��'�cف!K=���	�ox]�C���:���CƋ$�Q�EjS6�k�JUh=�o[~m>����O�{�2X?O�U5D=���3��͢g/�F�WҖ�̲�t�B��[��I��=����93�'��a�7� %�%b�ro��VR�v�����c�5-@�'B��P�z,��	������ϗ��m遫�p��#���LDI2��������cya��x�{^���� ~]5��^�1���.*��
/�5@��:���D�k�i*���(9�����^�kS�բw�G�� ��B�R�	j'�G�"	3��[��z�:��^�,r�u���� ��6q�}4���C�%�O�>�J7�櫕"�R���ަ1��::E0�(.>2��T�n��治p��$�6>.l��1Vd�,��?An��UE]* �L��e�[��@��]a�\*�MU=���	4=g�ne�N���"r���e���r����sJ"�UQ��1?-��U	�x!�P� ���K~-փ}�F�ӭ��V�cp�cTj6nN��A� lr��i�bXX�O�u�ּ�3�k��a,Y�5g���ߤ�{�Xύ'��Svv�/��28��[��&L���$TE��p����' �h�NJĦ��ސ��dՅ��?�*62�ڣ	Q9I�l�e��́�~�P�u�ޯ&fI�\M�c|�6�r�T���7��<�����E�l�f=$k��Wx�h�q�H4�ٙt2�b4j8<�L���q�գ�K!�m�b�Y������.���{�ʶQm�+����xN�-p+z�g"�G9eIL	Zmʔ'�e���ʬ��F5õ�J�W��S)��]�LA�е����쉫���5s�
�onj�eys�M��٫���y18���C�/�S;�o�?��xBF�e(�i� �`���-�hu�n�U%��Yp{�m����i��ʍ�� B!��BϞ�lV��r��h�z�}3=���ʏ� N�i[��(�����n�"���ƿ#��ׄ:��ײ�8nW܇!ӁP�Y�|�`���Nz�����9�B+���3����2W�(�q�btNE%�k�����U6�=.R���;
�����Y�Ce��{m.�$��n�j<�]���v�dm���P+�׷o�����%����%NW����7 [t��.��Q��:�#��i��V�H�#AUX��j�U����L�lV�F/r7'&J�B�n��z0{���3�N��� A	ol(0�55:�j%��!��5�a�X
�}��	@�h� q���2洀��(�Q��nFo��AkٝV���Y�؞X�����Fd�~ؑ�#����_�o�oiFi a�E�l�����=T�*��K�V��K� �#߰��;;H%��=՜i�gļ��i�2��4u�J��O�}��Õs�٠]A��w����d��v���W)-�����5J1Pz�:�j
�z����=)�5!7o*��̇��Ȏި�c�sQKnF�h>�T�!�i�-�[���&F�/�[L�;���Q��I5uԌ)�!]KZKA�ǽ��}���&��x(��;A����7�:R�^�d�*1�8ڣ�M�q{�`)Y͖�u*��)`����sp"�$|M�e8��YP��.i��b�Q�������h|͙	��P`L�'PXH�k����ΛG��y�ڰ5Ū?Q�S~��{vnj)�-_y�����e�ug�D�2ݿ>����@�h�E%Y�g菪��`�s���M�a�צʬ�i�:e4�`��{Vy���P�W���xk@��L����'1/���܃�W�%�!��2�¥"|�����m�]L�W�mQ����tΎ�ރɛG��Y����s'�k�� 6�R(��5�Xk�&�*�n�>�"O�XG���ܜ�F�|D%ƶ�V�)���i6y�V��D�ctO����h�3�]�t�)�}뙽t���-�%����_�K�����'�P�ս(E��,6�/�wr���,ad���]��ɢ�3oez�m\�$��F�f���A֢H����IG��Ƨ��b��O2�3��|_��O�����I�T����mQ�]��~�͇F�N��'���#�AX�懈XL��[N"bk$�[|�1��=3;`5x�"�2�8�e&�Z��
��v)n!��6s�g��+j{%Z�|k%������t܍�*�}`���\^~���d�M��Ƴ!~
�T�`�n����Ђx�34�t�i\��;�Ԋ-U"��NƼɣ��W̚��(��T�Y�{�#�P (���Z��W�6(nq\/��<#2~ �<ϓ?�}g�	Vs�
tp$5�[���O1����/̘e�^mx ěDK�?o	��	�/��G@��"�sk�7�/U{�nl�Y	��9����A�/��9Mp�J]	���[��l]����5?����D[�(C~��>/K�o�1��--�A�x,0m.��s_�����~���n-����*<��]W�%m?���_uD�<���91Gc�����؟��m��#����d	�~���9���E��R�m�Hnao4t�@|8�hm�$�Az��rp,qE��mQf!P��,�$�f("#VD���U���q��b�kf�H�>]�����!�p����,������m��l�����.��M��	u�X]<��3�b�����R�gSOkQ���&K3�,aN�dC�"�~G���r��tQx�Y�d&�|��g�Y͉�	R�!D�������N�К�|�10��Ԛc�D��o�f�xus1��s�8����õ�2}�<�
Qb$��q�h�YK�滅�4A���	��ݼ�h�磟ќ&�C�N��e'�����7$J��*U<M!���I�S=�	�`?>�}��"�	�`���P�������6�c�ÐW(�z������4L?t��r}=��ޑ@�O����|�.�0�F�`-�7ll(N��P�\Q���=f憤��P %��f�:�-����m�ۓ��/�b}Ӵ�$�?-�]<��k��s;� )/&�E��H���}�珰gm8��Y�F��T4�#�Ї/1s��ku��+|��4�C�ڌGJ�j;���I���t?,�����&ĺ�O��ҵ;0����F�/�n)��&����%��cx��{���8h�츢c���}����H�`�0^mT�Jl;iC{�6�ԝjk����4�Wm�]Ӳ1$ۥ��&De�Sd�ϳUO+�R�f�����U�u�Q�Rf���ƂY:�W�t�����{A�7®F�{�% S�\Q3�"H1��9��\��V�x������N@�j��A��7;���ٶd�g�?`�\ ���L��������Ȝ	���0�RN=!y�)c�ð㟃)v��)�ͷ���M!��,��%��6�9�H��1C�q V�ȕ���X�O�0��?*uF�nN��e��B<_;	F��s5���:�c�2�G��d~!'�(�ĵ�A�O7�3���`�>�i�p�fJ=�d��c$������m��d˕�kH��M�K��[Z���N�xS�k��2({ y7���|���*x�ml��;�*�8�/s����s�d�Ϗ�u��Re�	 �7P^+�_0E�����I�Is�2�8�_vŰ��.�Z�ޢR�'�Cr�J�v5M'�S>V�>k��g���9Eqo�y��̩°m{߲>l>�O�y~���6E}W����$��צ^������G��Y������%e2K����5��pz~WX�"4��7���::'bݘ�C�-%b����:���ș��{��5N��Z�H5�����n� �_ �
b��'��B@|$8�c��C��91���~�U㽔��)�����<�(E�7�\@u����o֥S���'V6  &mE�=�H��Hƈ����My(�o�A����yA�v<�L�������;ִAL�z%v��*ަa~KϞ�[2u�VT��;�9��Jj�G$����Br{&>e# e�y@�(�g(��9tP	f��������,���A:S�U�G�Ԛy�jAF����{Z�"��q��I��qi(��cd	�C6a�Rú�4O�U �c���ظ;�7V��$��L#���öB�% q�C|�;'�߼�ر@��"�vN���[2�������NЍA}��/w�������� �t�#)K�ٷ� y�Y^����#�'Q6���r�&�&v�(���W�K�{��&�ɫ�*�*9+�	`wN��s�B��̮Z`��Űq�b�%c8��r�,�\3qIҸ�]��X��%ޔ"r��W������)Vu��C�k��v6��nx�9Ύ���)R���1�s���@
q���5���wxƵT������B܈D���BwG��n�8��4�Aǒ�nu3�;	�fy;<?2cl"�2P�\�kw�86r�y��Q?HCƬ�bwor�?� 6��ve�57}9�yC*�U���7��O�{'����-���Ϥ��0�_=��+��;��a�?����@,�	�AH�d��ftj ��mJ�M�仡F�d�9��A��y3τ�r�{���o�7D�u0��G	d*����~�7t�H��ҵ�{�����$�C%��������F��
S�?l�D�IdH�)�{��R+��nn=B��ˁ`S�y,{�[�u���T����w�;��nӧe�5�j�/Q���[�?�x4c���n}Ɋs<ިW\��jg`��O)�ح��Uw4�W���ݫt�9H� �b�.�\��y���b�שS��
!���(��8|�Y2��ćf������`�jn��ט�K���aD�G�T��o.W4���s{��0�r�'QQb��i��t�t��� 1�b5R�Q~�i�X�������y`#J�K�"���=�t&����O8H����fs�i�a��*b��F�x��.8�n�X�~�/y]D�a��C \卿+X�o�z2PUT/�U<ݪs�;�e��D��\�EQd~5=`��&�6
�7�ϛ�N���&R7J�^6z�q8V�#r��9'�M�3ɁJM3W�?Oϻ����I<��,TL�����%X�B9	��
}�;{��<��⋻l�Ťo�Sm5~�YO��A@��y��)Ϝe�0ӏ�tl��n ��r�N Ζ!�K��.RJVo�=�l3L�z$Ԍ5�C��Bʈ�o;�#��m�!�%��i�x�yz�����<�M;x�C��c$�a�k��Q�Ap.?�V���#e��L}"�ض	�b�����E����Ů1�.���2���єR�b����;�lڪ��[	�Y����E-�]��(G�A+X���`�\"'pbc�\�sm��.\Q�E�O�E�}V���$�}�vѰ��y	���,V~��c9����)�?!�G숸K$�+=h�ް��R�g��C�K�_[�gRia�H��,c���4���A���W�D��M`-��SI��3N˷� �p0�(���+��դ$zta��R�?W�j���"چ=4��꧗���hy��i',I�\�I�,.�P4A�J��ԝ�� B
dy��?iY���N�v���ܜ���9�iКk��
+6+K]]@8�r%WF��MU_,�.���Y'�B�BQq����HW���z^���h���z����l��K���D����Dz
́v�E�v�;�S����a�V)6��rJ�ߜ�&���𨴃�u��ުl[�2���f�¦]�D�^� �g�?��:m�=$}0|���@���驀��=n�h2�=<�@�7�1����[���è1�2�v[K~�-�m�<?�N
ny�����m5��}~>4�1�#��I.��5���D(z=�i$�7���1O��f���Ӟ����%��b��%�3������F�$(ά|SX'��nl��g�X��
����z�}��Ya�>.[E�z�0JD��o��!��D�K�(<&I�'�������.� @T���@�<�z��D�P�C��F��q�r�FJ�6��N�¢�,T�o&�\)Ϊ8=��=]ڿ�'%P�w�<���`[�RK��rM֖<�׵d�ln�-_�)�<��7d5'^j�Pel��A��1p��*c���2q�9�x�Bs�Hfӈ��-D<�د)z�Pa8#��Y����!��Yw:9�Ob*
 ^v���*��Qd���E����,>�ZN�-h�څ�&�@m�t.Q2[��m��å�S+<���`��&^Wg��
�*KRN�Ӆ�Υ�ޞ@d#��os��n�'��bH��U�}��	C�4�E׋Z���~��-���B>ː��8=S8h��'�r@E%��*�L��;���e<M5�Lެ��oԕ��:���bY&po��A���]��ξd�&cE D�4D�&��b���R�s͑��my��]HdI��N��W���⸐�-خ�����|,�d[x�اKq9�7����b>z�5�e���컅>2\x���6�(y�~�@�Xrt�%H+`O�p"Tdq���׆q�����@r~��8�d0�'�g��|/eC����;���g�<>�K�M(ፔ�"���Էy���R:���5�\�֜PG��u��V�����&e�#�h�p�{���1��(��֡N��a�X&��[����m�QQ�yC�ߔ�C��Fl�t�L�Bf:�x9�_��с5��(!�k�ɂ�_j��L�V��Q@L�U�=�Ey����p��AQ�<F�ژ�.z�,�}27��Z(�ZM
�/C��g���UI��}u����
�Xh-��x	�����c�{�1(�e�� _5��q��n]"����u��g�n���î��!������V�"�2q���r�4� L=���N�,��.�"�}�s�������q�uɎl��WJ%�E�G��b<^P[��Q Z�V&���߲��pI�[��p�)6�����Y���4�?Z��ع̤��.�^����]������n��ҹ����5-���;�1�u���[7uF��;���Ez�m�e̓�X:�ĪnK����¿��GTq��y��I�`J�97�I6ɒY�;��<�-��lH�;�U��l�G
�r5V����da��o9��d<1h�=r���[D%��Si:��P[�o%��@�<B��XN-���y鵵s?b�n�Oѫw���iz���M����n�$��n�U2��(�'�ܽ)�ֳ8�0������V39����J�q�#�<�z��l6�f�)
W�EY�#�v�.Z�nƙ2�z� ā}��</�m��'%��i���+�d�����)=i�_�B{}t�moCU�`��h����kh��x^+�bA�-��o#�
2��O�?�z!D�b���7��s]�RxE�;�`�ƨ��`���!n�1Q2�4�ҽ�pF-�=������Þ�H��ω��ĝY�",��$��P�F�x"Kۊ��sL&J�d�;W��l��+���3�c���X�G)0&��vH���e3~R�d����0\�.n�H��ٞ}����X)�}]]���@���2M����Pwief����&1yF���La��+��W�O	�]S�@�K���:�;� �J��}���}D���J�(l�썫,��>��\�r�&��L��=L�!������ԇ�=(�s,���X�r/��� KR�J��&b�/MBP	��1/��j�"�A�ȕx}},�>�;Z���pc6E�o�����3�=�q����9��!��K<tGGa#�nW,<`/���P��D��
x��E>q�ԩ���uT ���uz�c��F���h�I$qUӵ��|���iZ�]fÕ2���=B��)�\�GK�b����u�c�;T9���V����xݾT���9Imt!4c�m*8/����𚙍,�\'�+���b��m�
Mp9�̜���Ԟ�ҩn)L��l�����7}Fc��z�'|𔠛��B��S<�6��G"r��r���3�͟���0�[i�:O!�; fO"߫�9oa��А�,��qG�o\q�N��h�%�i���~��bC8Ri.y\�E��wޖ"4��V��'˴<��kPRvb&��5G�]���ݾ�s����4�|S���R?
�"L��|_�)T� K!�JO�	]���F��>��P/����
ڥ�p�M�	��r8�N�����k���1}���~C��̘}�MW�w�����y�1�Z�N�]TH ��j����"�r�t~t�����_�JI��Z_��5-m�*��	���˻
فiVv��h|��(;�knN��S���5ý�C�w��������'r����z��s�U�I��#E02�\�L�:r��J-��7�?����3�he[�ǵ�s�B4���$C�Z�%�f���W.Jɗ�ܺa���z:��lU�n��ŋ+��7 [49��&7%�x�������l��`�&�:�j�E�O�#�7h�+����?;��AY-XOL_dU��L/��"V��"�_q�?Ճ��6ڒ[���g��[����=I�y��炍�$����B�����n�w*D�����-YGZݲC�����>���h^���4��P�#��^p�Ϛ�U2�O��!E�� /5��8jei�ѻO=T�Kd�����c��DRi�8�~��W�� -BH �S��@�P	�Mv8>����R����FJ���fhV�m��NY�Z�%���HB�7�Ԣ�v�s�}k�6�@�76w�#��3���;�����B���2�f� ����.��{˚ ��
���hL��b�I��8 " Ap�ډh�J��BZ�T��2e�k/���]VR����`����cY�T! ���)���^�z3z� ��k���E�����1v�kD��<�3|��q�#[��Oi��z<0>ܪK����_�
,v5���M�.����ʘ��bU/�ʻ��4�=�	� �c. q��Ǯ�4�1-c����q�URK�c+���Jw�L�ܢ+	vɉ�Yo?���=�!�c�
Tdgo'�Q[�~�o/�B����-�e6ꕪӳ� F&�8�6������e���$�{�XQ�6%��`Pm���?S��;��wՅ�0�T���OA��1�� 5��D&X'�\%�Ic����:�~/��?���}2���@���o�b!����F�_�HO���2���ԧ�ǲ�f�n�Z�B��I�M֯v���3�CL���B�9��}Ǐ���eg��uZ Ċr7�	�{w�EA���l��Y�]��6�;�z*bT��e�	`_�����z��|gF������P���K�
Q�E�Hl<�mI��xl��=5�F�+��F���m�%h�Pk��T(��W���Ht�!������_����Í�����Z��!l��eR5ODLq"i0�������7E�%ƛ�TS)-GF��|(m�;�h/���|��D��Y����^��o!��+�V^��k�s����(˹�����@\<g����򠞅Q�I'�g|ڒJ�}@�l�E�	�X�.��81������Xh��~S�W�r��{oPU{!�"z-ҝ R��v���qV"7������R�O��U/�x\�r(s���OCW��_
��m�vS�D����b'lbԽ.]�pW�6K����R\r�q&����	�b��+�ҼjU�v�*�1r�mhw�ɢ�;Y�B�2��4�:�N�e�	�լ������^>/�U�\ʗ1�E{k9�����k��\�����־׼\
�*�<�bSβ4�,��^�a���*�E/ _"7,%�v�1���t�c���Kx'������T�EԴǆ����Y�NuџH�n&��?EO�X��Hpr	���1��jB̀��`��&_fj( Ԋ�#�$O��o�`,�:��>?�}����oۂ��L�3�}:ȶP#����)�Y��­���ϘB$\ZD�\���u��P|������_��-_���f��	��7�v��,+�\~\.W5 /{ �;#���d�J�Cv�Y�[�J�?�������鞀t͛%���gV'"ZUz��x�k6?�<����_��"�zV*B�ΟJ��F�Wo�$�:��R�(Sk�?�5W�ER�c����(���L�O>z
,�TV�Xʂ��� �3IU�9��1W�h����;�NK*N�[��<4��l݂ҤO�,	��?H��U\�%K���'pݾ���P��N݊�+댽��I�!
����:	̴���癿�^�ʄi��E��L\)��C�g����"�8H�*xEEaD�f��&1�)�ѹ�=�.�8.c� �Z��mhp&�r���>	o�xc��-g��p�Q�i�2	n;�yV�Ve��S���Q��b�#�\C�;ὕJ������#��[U��@7J��E߇-չǽۥ�2��8{-N�l�Ē�+m��P?4#2������Y�Q���/��C�'��?G�DʪY��Su ��x`�������
����F���^�����k�@��948�zH�i!��*��K��a��.�Y���={{#`y�9��V-a��HEa�]?ɸw�C�z���;,p��!�5���`��+�vy�7��^��p��K>C>�����qc3�|D�R���,���ϻ��Q����ڭ���dJ��� ��Լ�n�����ߟr����E���G��I��0z�٨�����j�Y�@'�E��>�|��*��NŸ$��ub9�`��H��i�H�a[$V\d4 �WYq��� �
෱�VvȐ&7�.exr��W	��P�RLs�?G�����3�+���O2a��FG�,��,��{���u��>'��y)�w|����ZU��y��R7�����r�`�O�8�Kɒ�&�z�yl��g4���wԞ������g���>��.���V{kH��dO?!�@����j{ͩk�Y�B"D:����<�1h�C�z�xo6&�,�ٝf��  H��>\�wl"�%�Sq�5Cl���؄�%�����<��߃���-a���lΠ��x�H7b����R�hi^{ �X��r?\����ۡń�vŴI®�t;6�V��k�.4Ӕ������tcEA��z�Cߵ����#��y9	|��yG)U���N�D��`B��!2.\��tWmR���r�Ž�᧑`я&؏�/�M`e� ��.k��Q ���E�㒅�k�>A��,r�/�7nz�mz0Q�oӍЌ�Lvr��p�@=�o���P��rF����Ȼo�jWKVT� /�G,�"&��.Dm���V	�i�E�Aow����w��C�0�#��gs��z ��SHE�O@O����z�K+��D���E��u�B�ߝ��tc}À� �ڊpv�(�Ͷ��/)�� ���K[Ϳ ���(��@u��n��Eb�~�1j%��8���y�Ü�C�k����W'��^\�@�v>Y�v mM:ig�(�n�1�8��VQ���� �w^��@^�9 �m�1�_��N ��=�_%�_	2��� e�l!B���Z�zK� ��t=�.'^�t��ٖ��_�~��� =��$�}\&��+V�PO�a�#[�S*b<<1)ͣ�̀*Y��l��B&<�x�/�1u9/��DTxT~8�uQ� Be�ɂz�Bָ��Inh]� ���m���͜�p��;���S MV_C��ܖ{v�6�(MP4��eZoY�����*2Bݲk�ä�����>B���e�!��J��>Z#{�w@�x�`��?HϾB������6[�~Fd�BD��=�֣���i�t�X�J�o`ȆJ}�6�lN+|�����Y��#%<>~l�g��,�0J�C`���0��Oj�؛�TEI�1j�	�c�t����+JIm�s�h���Ō�ۇ���[��q�NM-a ���ī5��Yh�2;Kg�>2,j=���yZ��W�.r�!��U��Uqh�K,�­uD�~��hr����_{@��|9RE,vw��� [�C�q<7E��-ꙮ�����Jz^CAq���k�'��#[��=D.�D!�>��Ek�G����?@^��%Ўr+��'�?��>��xw�ź^9���/�}�773�r�R@�K�â�����>	�>��F���KX7B��R�j���η���B��*��}��7i\P*�pfB$gmGQ� ̖�J�@��
�=�Y8$]�S����7�g$5
1�O,�����cꋖ�$�'J����AF�V��T�|a&�Vpl A"�԰��jf��E�C��{���X�7`�`�kQV��H�oI����������Z�ff�cOt��!>���[Z��j^�γ��y����XU$Ҕ,�pv�$����6���G�[�jOˣ�5^R� �ʡ�C�"�˪"���_D
_Ɍ��n&b
��U���n2�;_�n� ��N?�2�oF�I��0���ox:3����Q�D�����D����>t;����"����2*�tVQ���X��ێ�e����r�E_��#��n�!8�e�Z�Fhˇ�͢�ځ���Փ���.��$�Ryv?����r�P�d�����8�J�d��0sH�eOzj�j�x�0Y��'=� ǰiv�^���5�O�!�|L]}���E%��쭿�S-��_��DV�w��N���A.+�:����	�.�u�����>\�W�1a!U��>ԭ7${D?w���`�τ�&Y��%�(4߯���^.�#ޯ��	N�3|�d+:�nQ�őp�p9 X���c`�b��ɮ��6����~�H��[�-��-��EzF��Y�<��&%�U<���P�l^��|I+D��s��P��z�f#0
�Xl2W�k�:�sӞ.����2�6����V$��
k�C���2�a����fV�k5P��7���{�宐YfoA�b��]�~bx�ʞA0*��ZW�浍�0��Q�۽�m�J��z�ۮ)��!׉O�!��˃�c=(ae���8v5�!l�������ۛ�d���� ��ϸu6x��+е;��P�=�(�����R�k��y�>�1@5:Osqz%Rקh��b}t}��H��%B�}86��x��X1Ar�u5�s�b�K"e��ߔ���B	��&πج���� ʕ���q6��3�Y
���EVɷ���T:���AJ��c�~��ב
:��C����k�g�]���J+3t"���&�.6�u~��}���+ʀ��O�����/O�FA�+!J���=_G���A��J�l^:��nz�׎ELy�&(@���h�.�UZ)�v|�vnw�4��\A`��c��v;u\$<����5!�a�F�3����kփ�v�U��E�a�K���z2���}�#.i��zU����զSt�����^�j��&�&͝ċFv���kv��&( $s�6�XB���z�]�(Rb�e�f;�n�ɞ��I��,�	�i8�n)Py�!�N�ܴ�����������*?�.$C,�E�n!L�;#J�����t`�y�+�'��Z�,�97�%��Z�c�t¸5`'�b)E�s��T�S\�!���͍KO���0S�iڍ���avMAU�n5����wln'�\0���ǻ�q�ڋJ�%:3�u5�K����gW���AWQd�K��S�
���ۖSZ'maȀc�g��ү��Z>�0����o�SE/���6y㉣Q|==}�W�����w
������i<��C]��벫|�9���rޡ��"�k.g�a�Ұ�x@@�qT*y�,�?)���n"B���v;�ʀ����4W���8�I�.}W�d\4�&��jQ�\*g��7w��yh#8���� �Xc�҂�L o��2�0 M��ّ{( ��A����R(f��|�&�`T���H�2聖�}?h���]���%�@�W ���X|;�k��{�.����`��*4nǸ����L�`��3k�4F+��3�.��>�h��0�E����F2�J4 ��?��ھ���:�������@��e9�p8��8[�n�J��^�!/%.�񀦚�I��"�[5��3��(/�����d�k���i)����v�p�O�w+��ʢ0���d��n�	6)�v�5��G��J .a��
.Wo�5v������!M�UA����'�����M8� ��i:� qKW�ށK����I��p[�*�O=� 	4?V������G�j�ۥ�1[�%��ic������V~��ք�Pϕl���t�W58,-x{y)+v-4�-�Fo��&ok{�s���1����j�ʾh��b�|���j¼�d���X�h�K$+��[�d�r�
Y4�
k7��a��}܃�s$�c�/�K���n��r�
�Bw/�`T[}]##1n�~n��DlaA�>|�˦�_{��wzrO %#�a��OH��F�k�٣���.!^��{�����o<�1��k��Ga���م�>��ʄi�q���UIɹ�@���gUk`B*���Sb�����i�	��7<�bF�}���"}��ζ����-PtD���&�l�q�̫U�����;�|���%y/����g�8�$��BS�la���{?!&��*ݾ��I� >���]�;�����`"8�
4�Î(-{�"o�|��/H\�Ts�Hk��v�=$p"�Q����v����P:D ���QT���B���O�zS��
�:?��ӷ��OC�b�F�\F���Ӯ�Q?�]�c�� B�l&�y疫��c����H��Ԥ�y��t���޻*��͎��Ә���xu#�a\�H���;V�;�4�(w'; �v��k�q3i�Ja5��E
\t��1�d�����G���dnX�S��E�{�Çx T�C��K�s�WJ��7W?l���+\&�g:�N��h��Qc##ε�Q�V��F���w~��������X9�Ѵ��y|QDC�p z�Ak��CEc�N#��pM����2{iJ[�Q\��`C6u#ۻ��#��W�=��=�1��D�x^am�B�R�C5f��@C��`�U�1��Bd�u�Мv���̗��e�VY����-�xÃ��B�����qG:��^U)}ڴ� ��ie�D���ܾ�`�b�)J�&QĎ�����oQz[BԎ��_��5Za��3�C%��>��,�5f��eНB�/C�z����$��[�����1�	� �3�����oJ�����ׇ����9���ǈ��;Y�
��v��W&��[��3w�5����Ժs�+zt}�����z�����%����.�ú�t�`�,�샸9��/��<+΃$;�{4���dDF�3:̪x{X�C7[�y�ܜ�h�U����t
)Ӫ{IG���h��p@�/��O5��\I9������u��;���o�p�<��LR�m�jk䀗c���y4ۯ���&�uD��	9���$�~/����M����Iɰh��B>~bx���X/ �"f�������P/�.��~����s���+�S�ǐO�ǚ��s0]�Ei��Cx~�V�(Z�2VT�e�q���gDްٔ��A���$� N���ݻ�����Qa��թ���@�_Z2Q��~�Dd"3������そ����r������俔o<O��c��,���yS�H�iOf� �ϧ�����n��J�CWTߞQ>?U�iZ� ��e1�Ѭ�i��BP��h�w	�Pn��b�8_R�\ݽR�*  ��(>.'Lq��M�����w3J�`�KZ�p�H�`��S�G��Z$q�9>��֓ÑP֏.����ٿF��U@e:B6\z�^�7+]�ђ���%I9҂Q���y���
a'^n�)e�a9��Q���z}#y����H��N����穀����Z:]F��`���4���p>X&����q˞�ʹ>6���a��9~�q��z@Y(d���,R��UX(Bw����\}��yf�F�Ѐ(f� �̽�oM�1~/Y2f/�@�8�����c�� ���M���T���A���wNm�Xvov�^�3V]�6CxC-��(d����r�(�r�w5�d$���M��~<��Զ�����4�MFzn�&A��������oC��I� #�?0{َJ,Ͳ�J�Fj�Id՘��t��UT�> V*�x�}���4y@yLu=�G��]-��Of.�f\bu ��ۜ�����IZ��9��x�(i�2�@�s�����>Vf��uA��u��z����_JZ {~ez#rz^^6n�CG.KR'O�#������@��k׎A �gk6� ��
-e��H�~����PN8��:A����K�<�$�@E����)�萾U��%����M~��-v貿���.i��:��x�U�	�,$���� ;�2B�e�ʈy��(*9��埯`* ��^"�9����}�7ב�Y"������Z{�_!Ll`�M0I��~zSX�����q+Օ���k`L�P���� %�`"�<B�r���lg�Ǭ_sYYo�o&Wn����U�G'�]�퇵���[s��LI����M$� �!��1����lq��9}�K���.�
�ynfb�G��4H����9�vg��OeS�>��*=X�A���G�1k���6���y4fq�?�u�D�;�����:=�js��ĸ^���^n�Y����y�&@�gr��F>͋�$(>?�~:�w���Ro��Ǐ~el���p�D.����EVa4U�h of Թ�|/u{2�LV��+�0�|�-����X���a9�0��ڱ�|��zuA[���F�����0��K�KG�;=Qˏ�f</0߻Kn�`�� b �v\�@y�wך�(ޑk�̐y<��O�����5 �0v*���ּ'@,�(J�)��f${����� R�g3�;�3�H>����/���f�������a���[Y�x�X�Z r�q-vdo�f&c,'��}Ԧ��4� v$n<r�h s\yB@1.Ǉ�/#ZT�
�*=p��/�	�@�7�M�5m���҃���\`ůS ���������A;kp�%�8��^�Iu鑴�f�v�O���)�V�����4�Q����&�¨+T�c�u��澃2�f���䂢%�(:C���W���#C�eްZfξ(�J8�%�����,dȰg��~OD~PSN�!�@5ʤx�	��!?q[Wt���"�Sw��l��'C���㢿M�N~J3vd�3�����ҵߊps͆V⣓3�7m�h^Ѹػ�3��I�|򥿶r���p�@bw�?�AIW(����'���$jq�z��pn���_WTShSg�}e�MV� �CX{�P��k2��#lx��N�?X_�Ƶ�F$(��#����j�/{v2��a �^Y+��t�����~�9p�"q����:�EAߓ��ڧ7��*yD�	���n�+&�j�0�I��}#ۑ"��fv+g�ہp1t��ت��;P��)�b�a� U�T�Qɚ�	�YI���vg\��+NϤ� �/!�b19U�|�)�)~n��eܠ��@�ܽ6����6+#MP�8�Ig6���+?dFR�}�s��,ϒ�:4��	G�5� ��=��(�!���Ԓc�%rI��n��{������tiS�%�N���zn���kDׅT��q�,�`�6���rhH�i���ɡ��	�ob���?�c�W2��G?t����xc�T��L���aJ�s����_��I���<���в�H�/�8<{�[F:e��F�r�G~��4h'�*�A\�5*�"�(K��
a`/΁z��"�MOnWW��=��.=��}�c��3�9Ej�����]�V�̅����m^4*�~X�+� {���
��Ȫ�&Ҧ��x�����*�*����mh����	����J@e``_�
�,�n�B^��>)G�>=*~�
y��q5�!����we�ɥ
�@��6�f��b���������$1���4N��ϥl��O�ft�Qp}�� �F�/

�c&G�Cъ���t`N2-v���;�{�e{IPaTUcVT�A�vݷ.�����0�HʵR���a���.�]���c|��{�tq�e)�_l�0�h>��@�Y�؍��_]4��gn���^�8�ՏMǆ1�3��_!\��g~�獔<90/����l�TR>�ȡ���2�ɵ�4���ve]>�Fi�[��(����_���N��]I?��1,��vB����.�}��R��?�x�Q��t�T[hw�2��b��")�h�h�B�ߙB��F��ޟ�ӥ�˰T+Ctq��+:"l��K��\�s�[����x3g;(hq5�G��v�����E�8�jk����y�ڻ�& ��xh��E�\�ڈȰI�͊h��5L�so��������= f����r���������ti5g!8-�&=���9FϽߧ�{`V׎��0t|�D�_V@V'e��o�K�)SL?B^�ѥ�����6ފ�$�!�?���tBP�?4=�O��c*l*mxeR����'��wu�p������2�����UT�E#ۘ�J!�_�<u��44X[
9���D���F�I�=A M���`���Z���yEP��k�_���.X��5�@�_����z�dW��s=����
J�D�=�JX9J�?ol��N��#tAn���<�㟔�}�fäV���󂬠/T�O`Jzc�-��`�k�Q�y�@�\�Q�Z(��׆��u���㙑7��곒J6Q�\8����p��\΃��U39]�!�`��S��WX]��V�6�ix�]"q+���hz�6�?�{&�+��F���7����*��B���eX|{S
���ZvF����wBqsۑ߼�.p3��w��y�9���įI�
�% ]��䤽[�/a���X�m�5Ҿ}�L!ʂC@B��+KiX牥eL[���t��غ�O�&}���˘�:/�9޷C� L���n��ܔ⎇�<{���߻kf%%��?�#�=��O�1p�|����iTc)c=�E%#�o��Xb���}UJ
��b�d�w�Rb�f1:
�>����E&>���z�Ӂs*;>�G��#!�#�W��5����KO��P�c�g�\�IŸ ާXrU`s%}1�e�J�#���u� ��Bz��^g ɩ��\^K�5��,��ӆ\D횥�d��Z�}�E���#�U�X�7I~ѯ�3�я���_�B8w�K�S<|CS��ڧS,a~z|OBt���u���dFr�����Ƶ�!�fEy�0`G�ǔ��$pz�0���Gv��&�M����m	â���Q��wQ���"�LREJI�C�A�M.�dM�4&�籼r��߁�0h���W/��J&����5�t���f�	w�j�ઝ��\yO4�菍����7�oyz������*�v��2T�����x�Qxq�m'���`B��	8p��,"����7���S�bQ"p˵�X�'�]�ؤGtcD7**��r��uf�eCw?v"4g�Ƙ��ƴWZQ,�Ê�-���at��9jV|�>�K!+߀�����_@�rX;��n�9�B�M�.UA('ܘ���c�Ҏ;��EWp�������������Ys�#��)�P�$�k�9���:V_U���-P��Fhr?Ra�t�\@����\����m���!e�|7W`��	FLZt��>�-k��#oc�e�1�/��P���؄zщ3�Q9������=���G�P;���7K�(��i���ۅlFS�[{�Q�ύ=�U;f�sx?-x��o��
=+�Z�n^�F��o���#ZWN���.$;�~���&|�n����&�-�湋�.�L3�	��f��X��,��A��.���9�I�p�J����C����p~��?=�7a�ɝ��$����9��>���6[��kc���X�WJ�7�#�:~��u�T ��A��$�)�X"��`Zi&���oS�b���D�\��ǉ�uuר�α�>�y���Α�^��	��_�vC������^MN�Qy��QH��T-G)�Ŝԭ�в3o���R����bO�b��ު�=�~�	pG�����tү��K��Xze�!�O'���з�1~�>Ь�5��� 8R���#ȝ��j+oYpN���Όb��0�y�b�'S׿ �� U1}K�I7��g_;�-����Z���b҉9�ߍ��}>CI�.u����:�'��T?z��z%)վW�m�A����^�!9�>�<���T�@�y]��7�+���%Z�R8�C�t��R�c���"e1����9�J3z�
L��x�_	ΰ���^h4ՌҍV�яb���&�_��X���'���PD(o����F�O��: �vA =Of�	,���>�&g <](*���'[���!.�0����,���RK[̉���'=��F|�c=�3 a���B�-z��r���%SDn��)Z�H��}��yF�G��9���k>�v%l�y˛����d�3��pHB���8�p�aj��Kf\1S��ƿN�_W��]H��� h\�v)ҭ���y9��@ƿa�@Y���t��گ�"xM�Bw{�{��<IA��J���IO5]�ǩ�@�����wfc�a�>XۿX�o���hT�vU�"d��!��G� j��2���Q���{��۔���7y�'^� $a��n�^�<;P=�)����Ad�l����n�����8����'iV'�R+wj�F�^z�Lܻf�Fo@�Y��XNS��&�E)�~�
���K�M�� sj:�4�	�X��b���E���US��Q�.�1�"����&�ܚ��d|��0�R���7����^�r��u�"���W)��"5D�^W)
O�G<�6�	�O�ų�^б�p�����]���[���q��@��*�:O������}(�F?���S
)&.$�l8�LG��j;��Y����hIq��g���3�2(7}[��F���d�c4I5�+Sl!����:Px�^=їkwe�ء���+����)WR�%��y��(uI��|s죝�<��p|89W��ۣa�Y�==R�=1���ؓ&㻼�Q4G�Ǐ����N��v
�����&�3s�U��h[�)�M0��o�8Z?~��D]��Nv������K�B��Z�2*˅����Nog�<O�c�K4���d����ƂT���jK���Z�j-��YO��0̎_���S0*�{;��T!'b��홏>X@��L���Gn/���tP�V�E�|IcIر`�xd���}J9���k��i6U�O~ܲ��Xt����x�%�Q�:��H���!K�%��|1�M5~]�)PׁM|�>������`���Zf���Ð�j�e�Cc����$D�g` �/]-�Q.�n�1�E3�o�]Y�]X�F��O0����b��嚘�v�(�pة���s:���N������I��~���U��.97K[�+U;�|�w�o�^������@UU�?�����ַ��u#sIذe�7�{�n�˫9Y���~�M���H눵uʷM����v��v��)�sZNc��7�z��!�;:�"v�Ha�����l.��W��@�eJjRP�rg��G�?D�A���H�b��Z
'��>x>���*�*���;3��9mI��e�M��;��'`ر�HH���b�؄��@f��Ց��>뵰sV�B����5s����2�Z�����>�?2L��V�)� y��7B��c��t*o�5ʆ{5��_#^�o����ʟ	��G���)x����O��r��e��6���10e�0V�e�J�U�O�#Xu��qI�������N"�K�&���i���&�W�����Dq#�8#�l���5v�}�_���>uu^���L��~XV�~���N�P���i5���[�I����z���������!�L+�7
��.��e%��ڋl�YtLW�ׂ�q�������CYsz"�yaQ����Z���j��an�b�+Is|w+�Ȯ��o�k(2��{1��x	�D�f�b��
45�6�N�H�ıD�C��?`:�hta�6����d�Q�#�N��?��V��L(r��`Vg%�ԙX�&?���g���M͹i5ÒY� �������xq�Q��g�zЋ	���BR9=�+fM��q`�������Zv�EUq}�ںrET��YF��`í�ƪ�G'����j���\�3��>�	�?+䴧�����M���K|����c��-6�����P��X��KoV���p&JP-���cc��6���3Y�2�ɇ4Y늑f�6뻳p�T������O�|�k�c���A��UV� ؑ��$)������6�4��K�/�R�t*;��x��f!��,�Y*�@ʮZ��Y8�b���/��q-�7(-]����Ĳc��3�,�%?Xn���yI���/�kf�sl襦�E��c~�O(����1�5�3���-ý�N[������r�;��X�ъB$�#�0[�x�h��3#4O薿9��¤���z��{>�b�-Z@*m�p��gģ.��
li�R(�vvKG蛅��_c����r�*a�'Փw!P}$&Et|�(�j�>�	��-AϪ�_?ތ������~mN�6������L/$]�$�j�g�(!���8ܞU��a��x��;�&J��(�כ�:�j2a��81���s�qq��˹Pp^�S�K�`og�Rr|hu���_��jA.��/�e(~GL�;+*���goK(Jf�>�r�FSm��78'mb�pUq� �g�_����pq�yZҋ�h���^w�_m�z"Vu.�b��5�A�������u�i��yk��|���������?�JǠQ5�niV���>�e�/6�q�w띔Δqʈ���	�Oa�Yv��u��5��ms�z��)F1u����b{�q s��1Ձ�3P5,q]���=NX�j�e_���3�FlM`�p�c��-�l�����q�E��Sw�&v�6�QiB�=:O����侳�8�m��/3(J�xL5.�k�{�~�#���Q�s$���g���r�U��B�.;�d��@v�G� ��ޞ.GiKXQ<����Ⱟ��47���k����J���F3��t�K+?���oķ#F�G|���1a�;f��dFS#T��_����[��=s�.��Y��t��t7�]$���.��L�}�`��ִ�m��(�����0�֋dt�I0kJ���x	(m����1�N�a��j�]I�>z��HQ��Vo��	��^����vġ$��530��ے�vU���L�1^��j�}���^|��V��V��gw���4f� �|1���T~���ޒF�T�������a��a�U����^�%�4u~ ~ӥ���<ق�s6I���$�Y�-;�G_(J*�!o�jod}b����:Mg���N��%��v��pX�[��AX�1��h!E��ĐO�y��y�a����G�h��"��p�	^�S}�Nl�HjՋ��!7��?��ɜ�������Ǫ���0�}D���3��@('�ҥ�4)�#Y������T)@h�eNc8�4+jT�wdm�x�;qlx�K��x�����r�`'�Lh�� �����������Vl���؄�	/��pcնᱫ׸^pJu9�l�0��)X�=�Z6��Y��4�n>{�|�.�nf��ϐ���3��M�6���XjE�Z�깪n,�,)��UbI��C2k�[a���h�;�����ƹ��̝� s��t��!F�Ӽ��a�|�ʭ����1�{���C���2��=�ܼI`�Sp(H��/���:
��`�&9,�������b�6[A��I�$D�rv�W=GG�,ީN��tMI
��n���ѵj[}�H��|���鶿�8�캃��Z/�t��GI��Z�8O�1��8�d��������$����!HZb��s'��ˤRi@n��(��FK`ſ��8��?��޼�EO/�d�����w��$��~��a�eXg���d��@��سa0����U٫�#���Փi�~N�L�QL�jȬ��̾H�P��Zei�O�hJ{-3r9B�u|K����kZ�eP��w����zL1�@`R���=}d�xэ��5���;T��9֏�d.�J�U�H9����X�8y%��XY�;�QH)x�C?��k�TejQ[�DP6=}J#F̮�{����Y	��Y���C���s�l��)����M_�p�P]�X��J���GhC~?�d*���X�(Y��P��!c����l˝�۽Y�G^�#��NY�
b��g��3�w'Tfy��e�EԪ�,&p��e�Xe�ɔ��ݷ��40������P�.�M7j��6q�*q�t2	����D���6�����5�Ad�E2(ĜG���H��ɯ���â/��|��s��O�6�͛�Ac�l���
��I��M�N��9U��	~�bT��-�HP�Qq&7�(��lG���R��F?�r=}���fU�ϻ%�CA���`}� �(����BA�-J�fJ�K߽W�)xeŀ�_��z��;|�1�)����`c�Õ�ѶPɈ�>y--�^b����j�0'�2]�D�pEw�KD��Ξ��[�;rJ�O���1Q#/cJ҇�����n�^OP����դ��l\w��O�Yht�w���|W]ꠕ$5���16ҫ�'�X¼@'F��}�h���Og�hH������G8{3�]g���p���HE-U�)����=Et ?!Uc��/��B�~1}��$�j/���mJc~S���vs�+Gc�K�1g�I&��ͺ�1��aE����B��h�#W;W�)�3X��FB1k\q�"�nQA��6�d��]�Q,AxI�͒�hi�*���Y�E�=�	 ������T�4!N��)J�ɚ��w����C����zo�Q%x+=Z�ȫd ��Cm���l�p�N�7Uq�
<ᝮ�hS�$m�Ziz釲�)���ۋS-(��T)/#2r7.}����܍`5�^�+���'Ђ
�s+���!3�FP���Ϋ>R��%��PV-�g� j W?�QH�z�*�5U��5���Et�bzi1��1Xz��o߱��	wQ+z��W@,䜢X��@!��5���6bh�Ee)H�6�#GK�ջ5��R
����'5���q4)MK���}p_ګ0��^#q�aZ�mڧ|�����q�v�d1w��b����t�9'�W�`�6��(˽c�����\�r�޳�Ln���>}c��a��%�wic�bİL渞���箸���yNv�4���#�@�.�y��lY�{�
����ޣ~9����"|#�� ��{iHG���Ҵ���C�G۶4��'_wZ������$� Ca/��l�en�Fh5�uGX�Rz4.�+u�;��Pܲ�O~�R�7m�\�C(ksmI��G�vR�u��ۣk�L1�:k���P�� ��(�Z5����暖{w��F��WuNP�7�����thK����<�88>jd�}�7ϰ�U�2�3(IEZ��n� J���u��`{��AG�g9k��W�
5b�Y�({r%u�*W}����'����!�G�(��v��
uŔXN��EdVA\1{z����2���/�^	�j��t�i����W�DG���(���sy��YeN�g�A�B����.��s�x��ŋ��
� h�Ҩ��6��8�.So�Vݙ��]S���?��s�R��3�s{ɣ��� Ed�+��'`���]3�2ҩUV+1��C��dZ<чj����ƕJ��i.��^4����̶!8���J�R0#CYj*#Y�X�˾��_��aq�n�fJ�M�$y��.�'?��3��i�b�~�ѳ#�G=|��k��n0�� .(���^�Z�_C(�@ҫ}���k�C�s�h�{�ͭ�U�NdF���@�ͣ���ٮ�dӾa�,�(�(T���Έ�XLA�S��3y�3� fn����F������u�����v��r������>��A2�݌�3���v�и��h���V�p�B�P�e͍�cNxM���MC��t�ЯZN�q+�fi.O���nF�F4J1y׹�A�Uy��A����dM�n^�@m��v�I��F9�e�dI2kη�P
�լ���י������Y�N�?���C�,��xE�z��܊�[��E�A��(�6��x��B�>5`�~t�x��[|���[���`�U�~D�k���u�W5cAt�dӪhVK$�6~@s! N�S?W������e!hPdî�k���Rwb����`�%��mZ�MC����:�Bi�����,Z��ZM��}��Yb��W���?��+;}���k�j���Y����3Z�ZF��r�O7z�os�%��S"���lo���!�u{�,ۜ��{��F�i��1��p�3��k\_��>�����_6�lL�j���������^��vm���D����KM��:9��
��VL����ǘԤ�A�eF�=���J�����&M)���`�(e�Y|������������8���9G���%�C��UU�^ـ�,�0��ŖFm��b��v����w���#(	�=�ROQ-�A�s�QD^��b�<vof@ �`(�g��aA[���ā	J(]�����M5��?�˿�0̨�d���Ǻ
���S!�O�˗��V����i��{�4��8D4�@$/���k���v�7��B�]���`��s/pIh��/��@~�<8=D��'�7�
YW�泷�16ޒ��<3��C�hi@���֒���>���m� ��XL~��sjL=��ex�|���0c{�"���m){NѨHfN����*4#��ˋ��Z��}x2D-1�g�}�(�c�f����)A`�*��m��J/PEP9G��'�{M!�}[�����`*F��YQ?{��G(�%bE�,ϰ��N�3��������`��\~zzQ��#�x���.12��M�٬��RhA99��ې���\⬗}H"�U�[1��ϻ���n���Dg[ܮ��~�E"}�be�o��O��
�E@o�,��<�p���r�h�f���l>���8�4Xo3�j4������AP���pW�r�6ܲ�`�VB06'�ɍo]�Y�����O�v��~@�Q���~�N��7� �.�����:i5vgz��˝�p����4�R]v�q���"�?���ZC���Q�mǄ��(�I�s��q�O��x�VY�-8u�K�%� б	��4U��U4%E���	6*��
M��4R�Ľ���8��?{��m�5G��<ys(��N��D$ǻ/'��/:;?�M�� ��3��a�=�:+k��Q+�~h�͕E�Ξl�D��f�,��E�̨L@ �7��r 2�{U��:��w�ݮ��#�!�U���6\	�m��q2`՝� -,s�j���%n^��I�;���ۆr�S4����#�ir޳��9!�:��L�J�U3���WZ�_�n�GD	6�H�j=ח�5!�Y���v�T7El��HB��oĥ~�^�ui�����&A5Yq�*~8���F͕X3���=
:a�T8{}��2t,>�_�-5�;@�b��[V���ƈ>��z��lR$��B�s�A3� �D���t�j鬹�\�Ó��+�z�d5�����!�:hJIp�A�9"anh�8 �� � �N#�~,�e+�G�[���D��
�N����L2G��ۍR���GY�!D�!>�F)D�A��Gsv�g��&u�D�!���.�T��]��}���.!��/Z��"�{���W�	ЯWxio1\p
a��՟�]�'�`<�����	������Y����Y!mI�à�����V�q���}�${:�6�;�L�x
�븷�m5r{km10� �wm�6[q�"k[��� ����t��oW�[��%y���"�g�:�v�&��0�tK �c�-q�..�,� }��]G�A��@N��C��09l��w��7%�p~⽆^��(?��`]dMߊ�FL�2] ?Ǌ~O��M��7~OH�	1:,!Z1��#���# ��2�֊��ze�`�D�ݧBŐ�h=�Gn�SP��=!���m*Y�G���'kc���J'��@�	ZY�[a�|/���G�� /��G𳒑X�_��ۮ�?�"L�}�"ֆQ�w���g%4Բ]Gxm �ǽ���-���{�tf=vFF�JKF/*��f����I���0�:=ԅ�����l�Bc��;LȀ����^���3˿(D�>N�$��	�"51��ϐ��&4?˨�C�����C#e��p�~Q�"�Q�>2��᳻���6Q������:�FJ���T�'�����V̾���.�惁����lf�6�UE:�Mƫ���$�e������&2a�[�TFiڈf�Ŕ��Q�����"m��8���B$���i�^Œ�����?�lJkH��K��df�q����ͽ"��2.��	�J��B��b�m</f(���p���5�����|��q+��
/���+�y�KE
�L���q,]G��U�|�����!�l�W���`E�JU�O��,b����.eU�[�zg���H ;��m���e�n�q/�y:-��O|t�@4�g�\��zz�����O�v�)�������
�I���w���gNwIB�n�n��fqm�s̿�
�
�i#�
R��j\�������.�������"�t�.BZ�����-%6Ft��w)�p�ue�[r����i���L�P��+�yl�Q��'��_&O���Yl������%�	�2ɝ2t�����Lt;�	��*s�w�7�T�%��*� 9�@\�����r�2Χ�]�>�df�+b_Nxӊ�k#�(hAʠ�g�xɜ��\��jI��Y���z���֩G@n��=���WX�t3�ZPlͥ�VG�z$=@���������K�f��TC�z���2��	"{��rP-�c�Ҭ�7 դpS9 R�6��aZC	AT=m	�Ex�wI���{JU\k��fkh���W�
1�}%-eg�%����A(�6ґ7ǟ�?�V�������Y-jE����hȍ��ucl�W�1�6����i�w�,$X�cb�`^PG��)�Pt���Gc7E3J,8Sի�>�d~�%Dȉ J���O�7B���<���#��	gT8��}�����`a�Ox�(��w;��&���Oxv�G=핺�����l��<��^*@LU�\wu=8���c�!���"��S�9�� �����wU݌y����PK� ��%ߥ���y1�躞ߩ�6�ە�}w���܎����^������(@�~^��Bژ5!�Ɔ�lx%���@�/p=B��"q�r�JDU�!r�]��F�e1)A������h߃@��".`��>4�#�E����]p/�L�e.b̸ NQ���W��AHԩ��_Pa<R�-�H�������N!�?� � ���ətw�f��Z�]��	"�OMg�"�Bɬ�7����)��Q�:N_ewW�,~�gQ٨�#`w�T�!$�B�j|cA�3 $�۽�~KG(1�nQ2;v��n�j>���=�ղ"��*��ݧ����L�D��W���|����e��G��y[��oq�l���f�q��bjm�c�פ�q��nJS���9BW!4��}IBӹ=z�����A��ST�i�y%�ǧ�8��Q�p��U;2�E=��=�[�e���5�J��I�U�J�|^{ �Y�r��/u�2��s�<D��(�U���]YAA��Ɓ�hoڮXr��@��ւP���'�����K�-�b�k�i�!w*ߪ�����t��"#M� l|Z!�� ���o�CԆ�\O'�hq��K6g���N#g2*�Xة�P�����A�FNw_Ҩ�^���~|hd���Fo�t[��K�p�l�1\��)�	��.^SeٽW��]�B�e�y.�VX<I�r��e���W�h�p�	�*y��5/���u�@�B��*uV�L�,���Zl�J���0�R�t���B�׌����,"�#�����P��'���{ΈN�d��?�2?��`!dj�U����ht�5�Y�>;����L��L Ƃ�ug�T"YO�ِ�u��7`p�J�@J��L0��h�u͠S���PI���J)�������==h�U�l=\�{���G��`��M>�Hd����C�D^$(���Py���2G�L��><0o��f�,�%��wpj���=Uԧ����^�1H�D�C�Ww�
��T�	蛧)�Nf������z��r��X˹�'����N{��qϹ��v�&]A��(2��O�#���U��a��kek4еw�x��!cS��������\��zz��w)R*���I��l���{��	���m�{�/��_���xu��kk�ZP�m����N� ��#�\��t	�!S���������	�0e��N����E�&�N|��#MzS4�Y��)��_4�"z�i��ti�U ��a-��+
mĽ�U���4;f������J[�Ġ��眤~F�z�1���'Q�:Ā� �j�I�c���B�9jG��'C���f���A�Z�e	J��w��D�F�(3@��類{�t#��X�C1g�O�m�DO/�ڼ�%MG��OI=�a4ص������`�i,X	P�gl�]��}����9��MD��`����f..����#^����92ҕ��y��j��b���z3�KsW� `��#͖Ƞ�7�ʍ�0l�m!�����p��K��w�zf5�$�4�$(G
�/9��[����)F�	YX]��QRNf}�+>!�G�^��`���r
ԬS�r"���i�EL����y���r8���Ų��- J���;��D��wa$� �gl� ��	�\��0�n#c�cbAӹ�M(�ScH��E�/s��6g�����6e�?~�4�*ǐ����~7�U5����.f�]����U��L��6���c)��vG��T&��|f��q2uU�,���k�
ꊚ���gLŝ	#�hr5��)�N�U7D���#y�
1?� 2T����i�^MJ?#4��){�F!��֞�b{xHH	�D�� zeOZ��b�Q����d��6��[C�<my�By�/�q~����}-���E�o'd��������M
#ml��^nM��;��Jq�h��Ym��W�\@���25�7ܸ&�������s�i��a��=�L���=�����tF$3�ǿ��s	� :�>.�������4��i,�������2EG�%���|:��^lJiYY�*	$�D��ƹ��/�R	BX��|!Y�bj=*��Q�
�� =��C��c�bؼQZ3WK�Y�;��m��\/l0����E��g�
�MO��^>���?�T'D@7�%�r,O���n
R�,Y�����B����'Z���4A5>{n�#|]Y�Z��'��cȈ_id}�����|�+_9�y�!�O>z�N8���q�~Eھ*==xgJ��[0�����j���!�(�ȌU	4�D_�)Vl	ʚEF�}�w�a;���#��J��frof�۩�����>�>9�ʺߔe��u!A�5Bj�Q��/�d`[U�0&�j)/�h�E:���n)ݧA�V�����'Xf&�.�w{��eB��(�.n���]��N��<� �� �;�Tlt��R��ż��^��#�R���{���W�/�'���僟l@�*��º�7��3�&��Ey���'d�6�<Ҧ��u�_Wje8(��G9�I��ͱ�������YZU:5۝�?f�`�փ�h+JM����o��]�Z��Ѝ:�C�ɗ,ȥq�:8|�W��"8�$Av����8��ݟ��� c��
��P�NAr�mن�ɴ����A��;ۦ{u�q[��/l��q$�\�yb"=8��tY��1S~,r���4�A�U�I��z�;K�NУЮ�Z�f.�|�)6=�
.���h���֩��S��:.H�r4@u0ެd �y>��Jt8�L���MQ�u7��|������,��%�t�x�����e#�&�KU���.x�����Av#��� �mE��U�L-_���9��b� >����������E�T�5�	���7���<n�	��(0��F�j-g���4>~u�� h ~k������󯊢׽��E��Q�k�U����Ia�<�v1�"�	���uX��j��P*���
z9����7e�V�GQ��wfw����D�C=
��C����-���NJW
F�Q���0ي��/SU�lm	m�ɮ�Rb��rO{��%�9b& �Mބ��B]E�T�<�����y�q��92.���oV��'�
�^ɨ�T��D��9�����K+�j{.+_
Q���r���=[����ߛ�%+�Q�C�	��C��#+���:�'w����LX��q?�)~��|���yc�՚z�je���ɡ2�W{���s3��LD�Am;�+}��n}Y㴹dݽ̫24�@ L���� '�^ͧ���*��0))����0J�4�v7��}��Ĩ��Y���dO�!]�N����x͂�A��q3�;왡���D�u*����Hx>� \~�k��뾘���.&4v�%E���O?7��q�7~0�<�Ls�{hn�Wŷ�N��{m�����Z��}Ϧs����+ ��S��2FFby�%n9�������2�O�;�/��6K㺤UU��ѓHB�N��+�|�a��W��n�l�"	Is�;�`c��eG��4��o�X�@o#��x�B��SE S�[�����Z��R���l-EtSw�jBg��5�["c�B�^�"��n�R�ahl*����Hڃr�jq 90�Kܿ�����@����:��N���&��,�p~�d�2������5�ah�,L�Ī9|�8DŤ$���zW�B{�
�*u��F�"��?1�w�}� [[�n�l���(K3�q�j��k�qe8��O3;�;��@���b�`�j��+�م��D��g�e�q��-��#��.���h�Z�G6�3�ϱ�F21��R>hRp��iP�����n���<П��׭0�/��^�XD{1��ҟ�J��?!I:���Q����@�LCr�4����/�[^�-ʹ��k\��^G�ef��֤���J��A��h�uÖ7�������p�@��	���9["��������d�?�{K���ݹ��ct����M�S��������}3���R�TI����d�SNE3�6�m��>wcK�ף��0{�� $�c�N�K��h�����&���<��K���Wb��2�l@�n�b?�~R'sx��C{��������*׬��i�Ԍ-��Y�^*l��V��оl%�K\jv�r�(�c�&�{W�-0���v05G�(L�>}U�ԾJ��v`��x.���������n8B�<�w�2��ɟ �]�b���!e�������;��i�wN��w��\��F�A�i>J��_`K�Fg�0Y�G�HT�=pz5���"�?4{�l�ȷfI,fmت�僭�D/ױ��@�i	��)��t��fV�6���c����9��Kk62z�*���W 6�9P�-�Of��(V��:x��N���pD��Y�P��* +�� �A��Y+���El!�S����t�@_�ļ���>�����?����w�
��K�t*�j,IQHX�b�zb�cj�(����;���G2�u���K1 ���x U�P4��SK����9���)N���XN�P�\͵4dGnj�Ap����4�HtGnFn��:���4�ŧ֕
1���
(����p(��w�AT �`!�,:h�/�w�E�9(w%�"4��hNT7���rw1����<`i�vD ��|�H
�0j�F�_���K��J��=��R6	v�6�׽_������P�TD�j�9�*�^r��̓It��C� �����3�}��)���R���S��ݓӜ��~x�z�#:W��X�{ :Pc�]�"^�t�i�'�zD�c����CF!s��򗤚��e�Gھ���	6��Ѷ�Qn�i�y���ܡ��(M��
�Ð�WSý$�{��@�'��lc;P��یɧ
ۛ��+b�[SE\�C��~��̕��Z���\"h	=�L�+қ.��|�j�W���M�L��ݢ&��z� �E]@=�`�oC=Ĕ����7��K�K,6�c�;
ѧ+� ��h�s;��{�*s@���` Z/T`�ԣ�����cuEY�f���J)'T�VwUX�@1�<e 5^<A Ea�璆!_��7��4l����e���q��#>.E7|��K���^_���r�8n&���1_#�Ͼ��������`>��ɯ�'�`M���=u��{ϗK$�¸4ZU{��|�����2�WE�x��t���sE��9�?-P����U�xF����	G��S1�[���'*p��:� @�K�^�0:�
V��W�J�
}�[Y����]��%��h�bJ���/��7��ؓ��M���[K˞���E%k`!)�u����E���[�KP$5T���_xPDd��4�}9s��ȱ�<�&B#<�Bm2��fOG~Pv�J���8�C���yQE���	J�xp^K�v�~gн�+�K�D�	F�;�@9O�0*}�4g�e3��z�~�Z˖�d+���/���x���F�Q��&"�\��X�����L�i5��B�|W���y�b���$'�6YVLK/�w|/��dqV�HP�':7i�f�<X�`Y��J@~��K�Z�)
Y��� �y-��c�׆!��Y�P?~~��==�Ɵ����!��$X�2�"���<�������_��ѡ�j�$�?��6��v��y�gC�
�`Ħ�>!5��Chnl�b��%����$�_�	1_D.�	�J����h4�/AM� u�Qΐ���Q���ءd�����g�hR���C�Y<?�R��nǳ4�.[(Ҝl�8���@B(&��߳����tm����w	��g�.�PW�����[�r��OC�P��.ӣ,����d
�� 	�����إ9�*�p�N�cm5�M8+����`�y������Y+uZ��'Qg�3�~F��д��c+���R���`���W�J1Jl�M¹s0ӳ�H�OK�y�k�j�E"� ���MfT�Y��V	��fN���D~K_PG��!��A��GٖdD\��ol	���x�'�:Q��2��������\ee�Sƪv����U�KRȶ�y�����"�iUe�Z�aw9�>%��,�aߒ��|&�Ł��Li�\&�Ѥ����`�:o�EN�7Ը����**��۷�(8��p�8P��%ԍ����g-m���<�y�|�̣@~�Y9ʥ�:Q�v��S#��M��2H���G?�E���`�F0X��}�G�)$]Ф��ބ�
�f�g]e����x1����-�������E��I���%�7�2k��'��¹3�w�{d�4�
��>�r�Dt��~[���(S��J�
a h�c�:�� ��{� �UN�	Nia�.�����=z�clia����� ν�����6�"�A�`�_�ps5���D.p6�A��ۿ��45�CD��Lv��ɑ�J����{�{��)d�� �m�ms���B�(؊�W������jtgߛA��<k?G��[�}�ʞ�]�K)�Lj�)L�Vv�iq�����'� 	3�Ե���m�xK6!k�<�� /+ț�:�
-�ꇢ���n
?��*c��`��zV�h_�p��ʦ ݴXq������5)`~���ˁ]N�<�ք���%q��-
��INy�k�P$d5s��Nڂ��;w%�t��m�އ��'��q=���ޒ�@ڏU��<�(��	x��h�L�?���N,5��o�@�f��g٫�e�i���q/�o��:$o�eD��k��N��E�����:�)Y�̀.3�ީx�6�ˣ�6������J(LLX�I���3N���;�uȠ�$�-GXClY��u��([[������b�jq�-�-_&�g��M���yn��nK�鷺d)[ܙ22;6;�!�n2NO|�����`�P�xV�a&��ɋ���`"�8��'��!y�;�&$ZҾi�}��nZ쀿9T��D�7���b8 �P�N��X}J���8��S�/KhK]f!!�gBY*�1A�t/��Dm���pH�d�1��ګ������q�No:A��t�Yi8�>�m�n���`@  ����[9b�X�FRU��:ׄn���w���j/�1�(D��x����=_e����[�� �:��m���o�!j,�٭=�"��mC$zX���LpVyV;.��v�Y]��Njr^,rdT������{�3����Y�����m�5p���XY��%�l�J�k
v�:`�Y�o��Y�%@yG
�3TV��jK�k1xhs�I/�������B�b���'7ҡ�V����^f0�#�톑W�Ƣ�a��.Ϋ-��<��ʽ8��RW�U�CM؎��N����LJq+
�'�O��u0L>�/?�cē�\���{�ө�&���ڧ��9��/�s+2cyX�6�qQ�E�/�M �,�3�auƸо��w��8�=�p����A S~�h��w���
~ZC�ó���G�ٍe'6����2����cZ~�U��?�}?���i��5�
O�nmu���U��\���
��z�^�R�O�����.��7"U4�M���V�\�����d��:H��wi���������]��ߨ��сMh]3PIV�=����8.֔"g4����5!�3i���I���8(�#�[yؿ_Ԟ*�(B���Fd�QLx ]R�%<k|j��j�F-����5Y*z�@8GPr��U2Vd5ا"��\J&3�� 
�.oh�"ﲎ]����]°��Dp��膏���vWxہ_M����ou �Zz���倡��]��g���S�O"��!Z��!���m�0?�fU�>�6AM6�:���ç���o��|e1t>�
��MZ���t��〾��0�fe%��<�n��9�u�P�y���O]3�Mz;��zp��:�����1���k���I�]I�"�ފ�����l��^�_񤼤Z��g>��Q��F�gzTM��]�2���T�yWF�<�vwY�1(��MC\L�H��)7
���l�,�d�B���h�d`u*	T9@��Ī�Z��<Y�����dz;�d�$����8a�
���a1y�[P�8D�T����君��~��9JPz�I�U��GK~�b�d�l�ӡd���"Z�&�LU�(U��0�2�5��f9���g
�y�#u�#�����9����ʄ��4��_$A/7k���W����n��H��"�5cr�iߍa��11f�6\�"Zd6�ٷS~ݎK�]! ��4�)�`���.7@����Zt����=FEx����vQKVc�h園�w!s�� �2|��𰹫����}����1	���cGi<�oO.qcN���C�X���t®y����v�i�>��(�h*��JF�[��ٟwRX~�"�X�B��r�|N�b����]�T3�m�#%��wB���Pz�_9.�c <�E�L|�'�ٹ+�,V_��Qn�:O����Y"ޭ������[GH�+ʁ��\���(����|���3�J��ȢG��a������y��oq k��xS������l��"��uR���R��M社�����|�j�� (���¦dH�!���f�����w����#��n�	m�}�s��3�C�6��Z%\����0jR}��+9���a�믥��Oņ!7������?�	SB`������N�����:�˾�A&"�Y���Pe7��@�z�L,X�3~^r�SPC�{+�u��5J�wS Ue��?��jq]��@א#�,L`�S�9���i3�+~��T��ӛ�|�P9�!�z/�����HE�'��+s���Mq2d?%M��YՕ��WI$ٹl(Adx�b�(�zB�94Q[mp-P���|�m�:P4zҁO�8�	N(P�z��o����!�,5)u7���%�]�/*�?5-ߕˬ�jI[r�彡/U3qgy��_�X	�}N4�ڭdC&��5~zέ�GH�k�zN��e줲nn���G��e��],�
h�x:��� Pko�(8ƪ���u�{Y�QͅA�[�ŏ��P��h9�s�)cPZơ�y�(kJ�Z�x_���q��ѻ��%�����/JI��?7�a��v��.��bU{?��Y�2�w����G7����B�#����;����������7Rt?�mb.�W���Fգ>�`3�F^��B&&x��[a|B:%ĭ��/�b,H�{�qgJ���C�k�T�pͿ�x9�i�VÄ��5�萢�Q%���  g}t�=�@���Ų7��=�G;��a�����,�,0��wZ�-
�,2�4�ki+~䗎~��v5���M���HU��,ERk�R"z�~0;�ϺW�gw��N�=����]A�E�&q72!/v+t�3�b6L��")��8��$s���w�<<�*{���VT�R�jW��O��3OU���?/-�	xt$�'���1��5��?�5T8``=p�=�����|��0�amB��պkB�f'#k8ɕ�!=FqOiq6�&HYù���7����^��k۠�����_�K��^2�,�)�O;�Iz��.�a�z�?���6�$RY!�Q��2��~�	�K�#�>��s����[ʥ��e�:.T�w)c�UP�G
h��U�9�E�E���B-l�_AZG��� Q���tM�g�>�����U����ז�T��N�\�w�)ߘe�){j�_��r��I׹���O���4��.�06g@�DP�׺=��;	epU�����`�J�Pjr5��2��I���R����`��]��`\fԱ�����\iH� D� ����eл-Ep�Y�Mm��ʝ���i�j�����Pr*䛰�&�,͢2P�/����Ĉ�砻�kd�U�AFo�,|}�O�`���6Cr�2�K�I�>�#�pR���5>N����(si9��8m�Y�0�4� &j�N�[a7��KۜU�˖B��`V����Q�����6ﺧ�7�R�N�?$X%9����*U��W&�w6
�i��ڽ;�M�	�^�s���qel���o��\B���&�$���TX5�����(�*b��1�%ͣs�uЄ	{D�8-��
]ť8@Ⱦ9y��ڻm~e5/?G�7�H >P��<�A�Og�ƴ�3{UX�a �������/�����b<�/�n�U����$����W������A�ON*���V�긡���V�5�=Xjj�ϻ�>�n��\�S����0ZĊ�H:�jl�zU�<��
�^�0��*rV��͒�hg�u���Q�4����oz(��"��dnl-�@R"�|N�%Q�9r@�c�X�����ׁ8/��tn��dY� Y�L��z�����4����0�q���ձ!x��Kg���ZER���y�&�ޓw�O}��-�P`�)M�
u���-�BTd$<@�O�[�n�z����"��"	f�R(�{K���R,ףd�Zbdr5��2]T��M�����ZFR��]�:O`�9x�~�L���.@�*�ֳ�۲u�`�*����Y���.&��E�n`�1k��0竤DDL�V��l�O]��j�lm��Vޏ��ӑ�eR�c#��Im���'T�~�թ����z��&�65���N,cr��l?.٭�4��o���B�"�g!���c�bQ����k�>EXc��՚{��x��ᒀ��^k�u�����u�b�V��t�ї�.��7��X�8�j�A����B(�L���( ��[W%����Q�V_R���om�F���_���&���c�@v�d$%9���9�l)�
_��	d�K��V���]��&['��x�[$���<suj7�����>Uk�q���߻:�A�〶��ڃ�&�Q�S�Wj{��ь=��-�j�TA2E�=q��u����P����o�@h�B^�G+Avݯ��\ 1�S�Y��R�7�O�y� V�J�	(��/<�٫�_����+WW���e<˟�Ov. ������A��A���]ę�k3�*�;C�ɭ9�i_���yv�w�p|(t�3~����2� "kate����!� �7GH	1��'#:Q�� m�R��Q�Z^� ����~SYE�R�-��*���(T�G��ܞF���˳��}��)��^`��
4w:�B���dd�3�۾ .
�����D{_V;�ALս(��-�f�V���k����	ʚ�(a=߱T�[L��jug� � �"��$\[ ա(J2���~Z�{�� [�|�l�.͔�ñ��f����E��j�(`Ɔ�cţ�I�� �ǦP����H��5�F�H�8�!���o����͋j��U+k~Lr
�ܶ	�뫐�~\
��W�����:D�f*F�1�\Mx��c5+g�Xʙ��˂1�55�  ����a;�$��]ԋi������%G�?�k�Зg�lh��
0���}�ד
�c��ګR�/�Hq��AF���k���{���w�OCP�zS��BS�+�DK�v祟\��LO)k�4^�*����)���ƈ� B}�Ncp{Hw�q9l��
/P�Շ�t�d9�mF�߱Hc[�\�� \R���n�kv�<%���F��D�A�3	USAܦG��ߤ*:\�"��2�8�S/�ܱw`�������l�(�umݽg�B�Y('
|W=U�1TK�l�n��������z�aeky�����}@��6�?VlIR!�pY�,�#��f�1�Y �{a�f�T�)��h
▪��.��� �S�K�g<��~�"m5.Y�+��f$�܈+�5E(BIS"�+B[!ĥq�h	�cKr�2�G�)�o�l�	:�����ۄ��A.�\��jO�܈_3��x��X���lT���������)$��d��v����@cv�X�Zf)�ǯ�y|��<墛Pj,Jb
K�}ш01Q���B�?y�~ԷL�>���#�<�t�����VR6p��Mf����c�:4��.�G��6��(�t�nM�����ݿf5NW�w;�"� i}ϭW�4�[��6z�/�z�w��@���dFA&�BkI>F)�~�,�����ҝ
:�ԯS��ү>F}�*�x�?�a�54�_'\#����n�!���iY���G�z�% �m��xv �|��P����>T���\�� �y٦6T�c@d2GำtI��߇��}�?���ݤ��#�>''y$���L�7J*�E�s�ʥvIז;�[�owcӟ�#��`�ǂ��q���J���'����,u��h���-�F�V[��`Ф����!�6b�f{p��뙋rS��� ��3�%�F�};�p�耤V�&�����Vw��U�J���8U���};R���t�f�k��8?8O��w<�B��1c��A+��@�?�dx ϩȐ�`��_�\�R�+][%0�/V.�}�2Ӥ��Fۆ��l�u�	-�d@!w0���L�����Q��Ǿjû�x>BWk[B��"����b�L������/Q���g ���,n���	$Sl��G1p��a�'�P���۰��5�W�^��K����;x�S,��#D��7o��r:D� �a�>HӞ�d9������E��g�v0$�ZMM�� p3^����[������߅�m&I*������s����p:p�"3V$�#`0V5$5�uߦ����Ο�V>��È��l�h�P�x�W4��*ZIOMC��@���7��Q�4Kѳ�����՟��(6����Tz�X5�]^b^�Qd�'���hN��`�
д?/���T�9��q�$]DM*�g��Hس�k[)����Rb�)�������7�?v�G?8��@�)OU%!��h��/D,���KV��2Fn*�d9��9�e
d�m"|Ĝu�N��b���p����/� ��c0<�X�y�7�A��OSo�0��1��ӰȮۘ �<�&��p嬶x���c�|� �葬��	�$+d�l��'�8{C�7��b\T�O��K|����	�h�n�����U+��U�V�u���b5u��1l�UP�X�Ry�p�wۑ���)I�w<CH��A�'7e�%!����L�����|�$���4�A����{���ﮣ')��ʯ��fB�8h"�����#� ����Mớvڞ�n�N��X�$�尐!�,\��i���X#% ��a!����.���^KʧX*3���}lf�~�C�Ʋ�0�I�T��R�"��EY���x�B`�� L{UAr��P�Ȓ�u|���RNԍ �@���	h�2�� �MTF�J� T�oI?��˺%Q�E�)'pBWG���|LMU�x[o9 ����ϵ$����Vg	�z�Ǉv]��+c�z�+sJ��?W얳Q��cd����L��z~H��xP��Jmد�,L�K�o�[��xW[�dLq2��?
~�t-,,����]�߅+�S�8i��+^�+�]�&��Q5C�N��ɨ��GZ?}(�X�����X�R��ϡ��J��Ε��hdN�1�5��_�z������Roy5/6V�'ʹ�����o��VP#�UaO��z�Xx��HIx��M|>@�����O�����}-��2�H�;5EQ��ë��S��w�pIW%��Ĭj%�������m�G��\nfFQP]z;E�ʢ�4���H ���&�>��i�m~:1�-�W8�����o��k�Lt�B��?M�{��,AY��_3U3��0̗��D�Nt����nӋj�~u�v�@�2���l3�����ΓƱ�e�-�k1{��3�9���Pz�����7��p�]�*�c=���o��i��^�߫������E�L���Q���$v�\�xWM����p�ƞz�LP|���'�'RJ&Յ�sE��Y�((5��f-�~�����96�c�F_�̬U�Tr�#�l�G�SWD�>`K!mhӾ:���)h���Ա	�O@�P�A�d�N��wFiJ�߶P��y6�w����/����tj����o����Z'���i&`��^F{���q6���~����r��L��v�(��9!����gEg���7���i4�Y�n5æ����D���ύ%W�t��Ϲ�Gc->��������X2�:�LC��p�N�y�����"~�<<lI/;�����n�=y� ���e*h 팥~)�.������"R�����G$�yLȐ,y"j|�X]l)�U�����D����0q1:7$�գ���@�.��0k�#[��5O̟PV���L�c��0k���!��ɫ3��m=H>f�0���BY##��1��H*y����W:\���t0~��IqY�d����B�JD�06��p�E���8�%P�Uo8�>�嫕wg��r�,��1�k��v؀0�bH�'�O.����H!���nR{�2�{=����N�K]h���v����
����������;�߀wW[B#'���>�QgiD��96K���or�XG�ҽ�cV���<�o����f��'��kM�[��`Y�$�œ�q�X��yz��5_�e�7 	��6P�F*.�S0�c �`TR����i`�-!�����Z8�[L���R~lm`��������'���
2���L���j���3���0�uq����u@��-"��U�q�}@�'ͽ:�Y��k�@p�R�u��@���_ȴ�)Ɵ��)}\�葊�4D�-;�5K��æŁ��Xnl����Gs�Z���+�Y�1��z��h�D����#Z��Kf���?q��IZ'
�hcF�fZGG�����(���G�rsjr�Kԩ7�(��� ��bW�����/���û�(i��b�VD��8���:��6ve�����	��U2V�䖦w�=���V����xZx5.�B�k_�+�M�s]0h��YS0�����sg!vc���jjN:��G�O�&�F{���]09�B�����b�G��C��̅�͡<�� �����0�*x�X� ��I��8!�ҿ�=�"��s��p�i�Z=��E"N[o5�E*2�'���� �CL- ���9��,�+繥O8��RӨ��!?u�����л[�Ǯ���N���'��x��q�	{�0��q#LG�?�[�ɾ+>�g�$�#,x�k�y�t;��ޞٍ�\�CH֐z�� ˬz脎�*_��!���"1{�"�_Y8���n`.KQ���5cf����]�;!�>m�v!R7�5��^,�>+�Ƞ ӴީwK	����:r���y.q�8�֣��q�n��5�$��"��I�
ݼL�!�J	,�JA�<�YV�ⳗ��W�i}i�ϰ�vk��q�ce[�R�Jj��zR>������sԂ��`��@?և��=��I%����Γ^�J*eQ�{ׂ��{�S�( �T��0#O��ћ��v���q��A��/�w e��dU�8uT|�����
W&��
v(Xy�䙎R�V�?�LiP�'岘{����u�?zTm�uNI����	U}BK�w�=��;�엵�E���t�%���Q��FceV��X�@&���(vO;h��c�įeQa���gۋ{k��,��1����(&d���^*��=v��<d1D/6S��9��P�������^>�x.�yt"�V +�!-s�'���9�~�T���<���������� 1#V�����P�~ۈ�!����}�/�N
m�v�;W�����Եo�)v�����;��>qͮM��,�?"�6s��9(kͲ�v���fJ"7���P���1���2C��C��Ɗ+y��"�h�ky�=��Jd�y>Thh ���|q}���l����i�+�����x�ev|�xȀcd�3 8���ʘS��>!���L��f� @6?:lHQ���k�Q}H���+��cNm���@j�U�ND��s������Ü1�䪶
�{@$���5�O����E���"����"��p�ʫ��+)c��8^\��co�ͩ2K��5�Ú���"�F�OdO��-^Nr��+����/�V� ˍg'��at���#� ��vx��14Ў��|R4Ns�n��Ô���]��Hp
�.�	�	"��fS��Y/J��N�bh#g{˟��E�|aX v���S�C�hoBm8�aTn���h��@�,�g�M����0ޣ�#3�T��>A�%�Iɔٙ�58kD��#�4J%�f ��x�3����4�UK��nJ��F��-�� �t��/S^8�Vl�������$��V[�|W���C	����Ί�5�,��%߭s!�1��3޲t	�0��W�;���5𹀈L�������/EF�̮6j�酸8KQ,ld'NW%���5*F��"����}�� l�>��'f���dA�oI<�����5^�3����4�4Xgg\���_]�m�ݝ�9�e���W���2���.���̣r�.�~�Fc�(�X��rV��qj�gz����Y�Av ϡɏ�o�R��rG�*�l�<.���"��R��:H�8j���&h7d�yo���9�QR�{ka��$l��`�;�V:iN����y�'w�൛��ј�W�Ub��|vW��k�XL|���wo�sJ���'��u�B;A@��x������Ƭ#��i,�@�G<���d�e��������E.k�� ��r����X	��}�Rs89�f�TJ�[0T?>�i23}s�R#�y�e|�.(��kB��d�p��:!-����Y����V�a&a`z������HV��|�=���R󞶰�7k�!.��g|�X�K[s���Xu�����N�U���#�&���Xg�a�F�ĺ��t��M���ݔ��>�l*���|���I���đ����C��[�fK��>{�u�j�z�dw��u|^��L%��5`��%nG}���\Ir�@D�'��l�WR棱���c�%�r�t���L���Ukv�r�*��<���������`����H���V� d�|)Dĉ��m��Ȗ< 
d�@=at�B6jY!��'Ol���
-S�����}j9�=�%O�7��I~I�BJ��!��3	fX���÷�Ի��,J�r�=��wa��a�m�+���%�R��&�jj�?@4Ռn�\��g����#���2�ɿǊ��䪑"Z�s�w�mg�����6����7/hUT��:�K#����؃^�����4�0v$���W�8@��ag� <F��(���J=�9���Α?�+��fb���%_��[_" ��J8.�筣��5HS"Q��\m�=J3N��G|sM����Aw�t&�5�T�t<B��2��cx��ꢨ/|!���}T�����������߳��[\�(���$�N��~F�������h� 6����m��Wpf:�c \��ǤG���"H^�>H�ª=} ����n�<	6�ݱ=���B��(q?'xk�]��2`���d]�3���������_���|�B�
/��yO��oh����F�������c��-�9���ai��3�4�[�����D�%���cCc��� ��ME&��-k9;�L�,���X!����t�H=>��v��N��~�L�s��Bdfج��]��w��S��^/ Fb�����g#H��:��7Y*�L�����&�R(D!�?��(h2	��������� ��nl���]0B]��X����Ŝ��ɉ��Q�T�P\�� ��Iq-�:H8JMm{2�:
�'U�	�ڧ�]����*D�ͯH_�HΜ:��gT�Ǣ�&&r��;k��Q�Ԗ(�֘h�Z�ѱOk����\��:���я��� �g�G��������e������>A�D�oCۿYݸ��{��M��l�1�����X�n�0���"c�ɃHS���]��0�M������< +��
䲟9
�'��l��?���L�\K����Z�~3��$9�<�
�免N�<�&�U|T!���lQ�VV��O��]טwM&#� x������������y�l2m;���2�WZo���0B|�h��z�����BP�� �x�{&s������w��;�n�5d <��gZ������4��~σ����,F|*n� ��V&$����`�8����&�=OA6?!� ����Tz����.��!|�������1]�WK1���x6�T��un!�ư�OB��<C5F��{�y�Y�^Z�/uR�w�l�p����`��_�E�4�i{�>�H'�TAH�����*���M4M�,B!2��l����8�x�I��'`1�4��<AX���&4��r���];V5�Cjp~߸X��ǽ��. e� �
;��Z0��<�p(z]��S�$<7��$4r��6��Ċ�k/��:���m c�S�x���PS�'�]�����4$R���q�g���r���xD��.��R��~а}F(A3�]�>�>�Ym ��1��J��T�Փ��_ 2izrv��Ӽ>y�hi*Tr�֔4�1s����1���"���ӛ�����]U���J��x�g��nx8�+�L�p�0g�D'�z��{$CA����5ƽQK���l�>�3]�����U����H�2���"�g�܃���Z��Q�@��u��[Z�.�IUQ1J,��Y��>,�> K8-��Y,~XlHy���U������d>5%�G���`F���H"�R�9��]v��jƽ�3�<�#T���c@p3�+��@�x�����5�|fa�8eR��[�t�y���C�T�/��g�U)`�q�Ox�skQM_xr�a3��$SP\�(��i��F*�)K�w�k�⬘�լ���2�z�2ڕFG�? '��u�����r�ͶRn�����X�$Q��7Iq������rh2!N,`a.���}�Mnѻ�m�?AQs���`���a������X�4'MQ����q2T)��y,�D�� ��#rcJ9T���.�����;��
(�U�<�e�L�\�PX�6i��'kC��:��3EP�˝\�<��o�5����$��⬞5(���@�y�����+fK�a<aD���\vkBpP�o
�Mx��/���?�W�Z6����/$sW
�w�b�\a�a����0��+��Ab�A�s�T�p��t���/�]Q7*^F�u�+}�~�<��T���ҊV=�(�~�71�j�]�1�RI�k�N�$@���l��^�� �ql��]}�U� Z�Bר~Ǒ"�[Uy�Hѹv?p5#׶ �<���C�?��b�G
�&����A���xa,i_@4�[�=B��F.�"��M$������։�(.�G/ˠ��K�1��4-�Ÿ�F�@�R���W,cj�x
�w*��e��ś@w�wG�Ie�Z"�����֓���0���p�6�����E�B��C����S�s�{��[e�������F�Yᔒ2n.n��z3�L?�����K>n&��-V�gE����<i�Yt:��s@���>���X�S��6�ߵ��sľ�/���Xy˵c8@���q���"�i6�`d#��/؞o˔ ������j�����ߐ�I��̏�mX-ז����ȏ���5)� ��u}ӸR����Y���a�*��<�"���6�w�v��a�}��[��Y�]6�out/�$��%��3i�����,�$>�)
J��,E��p4��(�V��+���=	�QT�<��W![Ɵ.=��[4~٦�{�����:eR%��ؽ0�<7�ڽF ��YF학u	;j���_[hp�o���i�����'�[Cw�c�@-*O�Ye�KM����1�U����s�}h�Wr��b�y��!�i~�y�}�dh�M���v2\N�m����i���<W�F.9/��7��4���zh>��
)�n��>����*H�� \'J���.���i,.m�{��'��s��r�My��\*���zM>������Q��&(W�E�w@�Fă_�%ޥ�Q.�>��Ͱߢ�Z7,T�Iu�IP�4#��*'�)_�K�r�^��b���F^���
A�=���K4+��_�F ��3P�iN�oX;)z���`�|�A����Z���B_PBM�#Ԕ{U�5n/ɩBR�"����� ]��nf��җL9'�ا�B%B^P�T�UegT6��_Rc�����G.h��h���ie���x�}>��D?����^�[��k��%8���±;qn���~�=Pd�t����)�$��k����L"P�soc7�egp��b�$0��B+� ��آ�K�QgǏi��4B���N3�O-�����H-E�Br��NG��UO[L�}�ܡ	m���� ?5�����~�Ǯ�h��w����|�f���$�Ԉ�3���b�
����KW��]f;S���_��T�Έ%�t'z�e5^�1��\�j�8��멜+�J�]4��H!�.�%;��G�p(Y�ȿ�Y�e�[;;hE���Uwl�}˸ș�tH�\�p�Zf��C5�v0F���Z�\�V��b�'a�_�@F�å$;��E[�������	!�ƭ]uO�ZH���au�4!�ֱhF�M��Ȋ��c�	�j���v��>�l8��B��ӎ��_�y5{�]Qm�N=��<9���S�!�Ȏ^ٓjJ� :���E������y���8�_��� Җ��n��F��6�+�uu��jb�5�9��מ�l҇�a��C�ɳ֠Cb��h���XF�W':;S�7Ah��������\��]g�/Q��3ь�'�(n�.��!�����$p���J*v(d�^;Fu1�|�y��1��6��ެ|�y?�M��\Cɬ�r#���η�R�CREM� y�z@w|�8�Ӆg���&��R��G"�X�N5%���_'��C��t�ĞQ�_�(?�`6q/�_eP.*��(D�ă�"��G�$��*���E�:�޶�]��+:��k$��h�iʛ��׫�����,'�	�NИ;J��ɝ�W_�´p�P���i�r�ۼzTj!=1%��g���ӊW8;O�w� 17����0�����}�=N)��/vX
 �Sl�"|��X@��:�zdϪ +%�>Pk�1]7�=�z�Qn�t�����a;^�n���������r_��g�,���g�.����K�{'� aoe�r��FoP��Ӎ�iC��p���j��et�-{v6�}ܱ��jذ������ܽ����ҁ1\���C�[��-|f�y�����N�_T�pNPz��CM��F����-�t]W��2	Yl���Vw@��S���;�.�����\�c(=}��g!M��m��W{�I<��j��o?��!ʕ#�2���;�:�O�?���w����zV���+:�|�Zz�ג���r�a�1vMI	�w�_
��0,/�7�$T;�F���gpQ"���^ք�l�rd���G�xkMT���\)��a ?C��bO�4Ǎ�[�8��%�M�����Y2��IzO������z�m�to>�/$�U#
����P��^D �==}�P���v��Xf
~ٌ#)۝�/�"	?�ȵO�o��&�Q�I���O6[��¨�Q����-\��8��;.��$��c|�t�4$��QO���fa����쥽+-}�s�GD9�Z�@f�����TTm������S@��J(_����K�k�KWR��`b��^�X��L�I�3���o/8�	����1�9�����C��2��/gY����%��5���#u*ܻ`�hbysT�۔Y�;��6�������X�-u��);�v#X�����wp�$ψɸ2�5=q���|�Zv8�m��ӧ�p�8�Z��1�O�+��d��l��[�q�B�7߬�$���*zˣlUbx���l7�YA�6CV#�އ,H��5W$hPW�R,�m@6I�!U��#A/��%�(}��ȵ���,�3bv�|���Y+v?��4���{T���� v���8�I� E�δH�"��1-��K�+��o���J��A��E&�,\*˝����6UTp�K��U��.�.^�� ¨?���4;���e��z)wL��	<A� �q�m�&� �&����7ff�r��[N�jg��)<�+x��-$��Wq*�B�f�� /.�k���.������M'�;aFc�ทnf�Uǵ��i �ָ�nQ6��џYi >���V�D�pEͪ.hr?���Q�܃�V���b|JG
��e�b�� rHȑ�]r���C3��]w�#,a�A���DB�%�R��b����Y�Sg��rB�A^x�)Xl5�R�������2��i?&����S#�.X�����ۡG)�J(i�r@�_�v���\x��*k�XU Qm�V�5qƀ"�������C!���I��*���*SK��b�����C��ɏ�!��$�2���?[N l���>��T��_�,ް�6��,x]��Q�>A�^���k��>�Z/�@��L��q�%e��+�u�3hÅ�z<�4�|�m����9�������[-�� ����� �ڵ)�$\�4���ˀ3{>�����]��i�g��?3���MD�~���~'CNyY�߫D/v1Q��f�b�������gE���ew��P�/�}��!u�I��(m2�K>�n ��5s	��e,�_�%�N;�_�v@{8B��)Y��d�������lZ�> 9#�[47�ϥȌ��˯_�L�Tՠ���őO��5��2(>���s7%���\�c�8(����� �\i�嶅Y�밒!����DW?�W�-	VT}c��(K[�
�WZP�-#M����>��M�&�M�=yn��_�3q:���*�In�)?��m���9���i˼���Mf��<�mq��>��)���C��/4U����%�\��]puw�ڝ.BG�EZ@�ͫ�E����t>� ^�	�����Zƣ��e���-�S=X���n�u�k|c�"Q?Cg1�X18��0we���Dл���
�~� wTו��VA�B���������P�3�C~�'AC'6m�{���F=��8sBV�: ���X{//��ܴu%S�e\f�ٝ��7cK��F��5;���guY��X�K����EuF�4��gI�pNm�vG%� �0��․�[��F��.$�RՐ�;�l|�:}m<)��T	(�$ b�l��)))H�d�Ҝd��K/ ПHe�5��<� KV������dŔm�N�����D��J�k��ܠ?rӀ��8q�hC�:+����m2Ϗ���c"j����C�VD��xH01(�􉴺���<7�w�6R�a/(�]Ú0=i;R�B�30�H��g�$O!(��z��®�!8>q� O]��I�N�n2=eU�'��\k����4���ku�)�5��H&��`08�ZG�z[�ˬ+�������	,��Pk���a�nŠ���ڿx��@_�e�d$�|���֟~c����r�`S����{�;�Sm�a⧼�-V�-m5TU�Q�3,��J�]��Ɍy��2�r�To��P�1�����h�`������	�Z���W7��L�N��O�I�="b_������r� �]YOO���|,�Sgbcnbd�!z�+����f	͛2�@��7+*�v����Z�w��^'�{\'x���^oq�$��lJX��D�E!�����Dw�DP�������޽9�߈�S�yP��ނI2���يj�B�Yvl0W[o���_b�s/���:�|ű0?�(+&�Pah:3�!��Hӕy�����=��,^�*x���,5я��QZE�]@L�ڍ�0?�LW�s� �W
IGϱ���ы_L�F��v'#il�%.�JfG�ml��*i�" `�R���^!�w��q��IW��6�<:Ou�m>����@���#��49��N&�|k,�q�yZCn��!��+�kiJ&�o�B��W)ǁ�����:�h�z"$�K�p��G��`�����i=}*Z�B�	t���!#������~�W�����
��R~�R4��� �X��ɗgA�ʈ-S��69+�Ч��7K�Tڑ��s*�$7Y�P�?�9�׎Q<���L�*�~����=Cl�Z�%�J{ ��:|'9ܽ+.�L.��{G�m���x(�VF�۳��2�ޱvS-�~�xځ|K>�tO�]LYh|'޻�*��m�� �p��K ��	�G	V�峖�%J�( \�+P����t�M��eʦ�5zBՄ�.R3�2�&ڑ�����ڇ��վe������7<M$2��{�h.	�p��\e�t/p��_���Z�y��tÂ�U�O��S}SLsD"�>����|�Ig�$Nj}'}QWW1*_��t�v�K��H�D� �B$�г0W���w��Մ<k��<U�X�l��4^D�\AfUL�.��zD��&�o�g�O�"�v��μ/=k4�����p�"�kc�6��-5d���;s�Ơ�jU?�؎m�W%�k2���}^7�ꫯF�Y��@�^�X��H�'lԏv;�:#�ύ%TÜD��/Z�U~��Ռ�bH��.�v^�bYۼ�+�p���6T2FJ����H���#V�c�ɨ�/��e�A��M��
��۾֌be_>���!3���r���o1
W���0����u��ޢ�U�ͮ��*�!�c�ܯ��;�.��E!E�I5��,ĸ/����bsm;]���o�HdA��"	?�)*3Z�%��T�&��~BRά��q�Rv�+0�>?E!N���`y��k�B�o�/O� ����6Y�ԣY_x8kf|U&�	�yn�B�񾨤=���T=wBvQٹ�AY�`��q�h=��_�S-܏�G���*�J^�N����Yʢ��((������Bs��I���o_��)}��!A^
Tp�\��\��vB6��aݚ����4�o.�Y��nH�I�F��[�{ ��a�H�rmwU=���^'�i�"�
S��fmU���-eJ}��2�X׭��F��7��l�@?:PP�/t��X׵��trwp�u܉�vCB1` Ql���Dɐ��T?ϭJx��9�|��|�_��pS7��6Ol:���>n�_��=E�(��T|��h�c<$��c<
�Y�r� �s����|U�:r�H���7V�&x7VU!��W��}�1*v���Z��`��24E<~1�*�s�dw���CO(C�=�j�f��M��Y���,;�޵��ܓ��N0'o�Ve���:��"�Z�(v���k- ��}��Ǎ�
i�h~!�޻2��!�ak�#~��X��yrn�?#8F�kc�J�̜�X�36�ߡ�HP�?��}��-�uj��gAPrXϦ��gb���nrG���q���;8���F��3&����)K8�`�� �,�z�*3���@��x5C�=��b�9D��n�R�M�a�kj�$ӯ�&���>~��JE��'�_�Y��H9���@��V�):���5^�M� �'�A�L���&�(w9���L�s<6����hr.��1K9?�^���7=bq!�q8��5x��[���ѩ���+�u�� �p�MP��@����=��1Q��P�z����J]�L��Bf�'{� 1w�R�N=�|��W����ά4ԹZ)&����D��٩�8wl��� `T�i$���B:��%Q���Mh�)�mR�y(f��4]D33
E��O���W�!gK��s��߹�Y��H���p޴Q�Iɖ�/
nQBI���yes |3��X?|�1���D������)İ�gYT��?���YF�c`�����y�B�?ƤP����}mB秕�>Ž�y�V�0�N�o=��'��eW�2�@&{�7�ф�P|�ky������	�ef1�ꥯ��Pҍ�6V�57S]<�lJP�X�xJN!Ƽ�*�j&$u�ׂ�>���daz�$��q��	͟���6O,�������,� ��n���d��ړ�k���ti�Q����IK�g��Q�C2%���m��(@5�M�שnš.c9M�4E��cNIF����މre/�N��M�/��-��؃!Y�&Cұ����M��9^�{ݿ�}�O6.N�_���3��jbKaҍ��|��^\�-"aaW�	J����y�N�D�A�j���_a[5 WU�({RÀBN�j̶k-�m'�7�� V���|��'�>ȯO0<O���sM�Dą���lG��h]�O
���V�9E��<�D3�˭02��������M����Y��7�э�L���րbh���F�g�J�mZ���G� ��y�]��xo����G1Z�_0�sn&:h�}3NJ�h�����O�9Ҥ"(�����u�+���r�6��_�k8s���ln�%��q۩P�������Q
Ӕ��c�	�0?^��j�u��g)��	!Ji]�y�%��(y8��^|z�E������ ���n�19n��\ƓA����%F�W?��I��9���٧���^�UK��+�#��r�g�v�U�h:6E�Є�Z�ϵ7{5���N��O�5�'�tN�O;(s�����M:ǻ�.�%��_=Nq�6�4>nJ���R�xt,����ύ#�{����>Ҕ9��s�ߪ<�<h#�V!��A6�i���E�V�;�����ʗ򊼠�5�mW�e�U��\!�؂'K_.����ݳn�}O�c����S��4�k%��}��{�33�ty%Z���)�����Z5[Gzu�R�����'�I$�9���9�y��WgY("��*����ۉ��wkY}Ӎձ��s�$�b�	�������1�A�xȭ�十&��
8tK�
8�I#�x��z�m_�š�yC���&=|��,�s�]�|���;K	���u�!�B~ 6ۗr�ܼ� �܎�6Z+q��0�D$��y�x=_Rk
����p�?DuW^�ek��j�׆���b����@���@?����L�rjM����\J�<��V{m���`�%����q#O�m�h��qȇ.��"sݰ5�TUh�1ѫY��e>�<�M�L(�TO�zi}aޣq3+�!\E� ==+nU�S��C�F��EkJ*�3"Q�"qϗ��	��������ً�j�#g�ZcK�p8]$��;��-�y6�{��M��ɗ�n��e������A�
�-���m4��vkL  �8���ۙ5�X��K!c�[y�Z��ͳ��
��`^5Q7���>��O��`a(�E����N�H/ݿ,��[xv�ǆ`��C�l@eU4N�����/0�'��l�tf%2X42��,�+��������H_����7�m��WYa.�~��r>����g ��1EE4��M&.	ʚ�#��/�[�j+�Ȍ"�}�
�&�g� f��ۛ��W����x��o %��j�?��%�N"�xZ���X�<e�:��CV���XS��ZO'$��:O���7�G��앸��wK�S,Dڑ~��EhLZ�Yd瞨�fS�Z%Dݝ���>m)����ͤ����bV�=��2](���W��NݫS�"�������eIT�j��T��bw� 砦d�����T��Ne���pC��?�-k���j4�L��Y2��h�3���E)^w���D@n3��>O��®�S6���I��󴚞�	���9&��`����[X
N���Ô�3�Q�ȅ,���+�]�#0�E}j�[�����V�.�{3bM� ]��xxz�y���	ҏ�T��!5�s�h�%�d�|R��#��{l�����ʐ�=;C��5�|#�/�x(���_��cVa׳&�YT����C!��tO.��u�,r
�^�S���X������0� &.���S)�u}�D�;F��U�B��ߒY���=�+<R�iu��G^���,Pj�ak�"ӵ���ql^�8T6�T
P:*ڐ�9;@����9ڎ!�G�O��qN3� HҔ���"��8��1����~q�Ӧ�ٰY)~r�����X�.c��=%�Y3kO�㤼�*��#�V��n>� �{cZ)���E����b2w��"�Ԑ[�TS�p��ɽ"���e��f�^ ��Y'�>ùpp�6r� ]�@y�0���E|ǫ:�;�=l�����ڢ��{��6UM�1m���b�a��۩A����2͠�����c��5޺��u�� F�-Ω�3X���y��)WC��4� ɷ�ȟ�lF�
��յ0�l���?؏�H5��*Y'��>M(D���ȦА`?����S��
k�>��\AB�	w���G�qix��Ղ��]���w�ɰJL����p���Zk�I�H�7�DO��%��D��[���k1�,���Ls�Ȓ�*!j�uΑ��
�w���I�!E/��I����܆c�~��8z[�C��h�u���|�y<���"��nH�kY0�ǁ�|�Z1�F)���]��o2��M`T:̱���r�]���������{f�-v���Mγ4s���ѪR�S($�H�����K�z�r�I�ck[�.�+��$S��^$eb�F8�g���zZ؛�W�f��?�!Q������l�˟�<�@%5/� o�y&83�;L(�׉�"�vέ漀�l�y.n�mo� �͝��1 |M�Њ���l�ŭ1��-��45w���Y|��f�g��m�_��lB@�P�><�&55h���T�k�UǺ���ꕝ�rp�� ƉT��R�r�s"Lr�{����㞲)m�Лq
{A!\��r<�Hc׊���ξU�m��� =��a�O�a�r9��iVDm� �P�/�vWe�DG��h�����:\��WG6(�І�3IT�)�Vw�zS33�~����'�W��9��q�����G���HQG�MR���Ɖl�{kħ�u���z{AȊ���[p���i�37wD��(�������j��g�婟x���,�L4%i\�+rfC^�f��b��t�o�H��A؎��_?�;���md���9UYD�nV��a�)A7��9Z�ɗT��|d�v��uF�n�sJ/�WO9oOo"�x���ܸ<��f˩�6��H]N̾)�!5*zǕ��\FQ#�6O��6w���u�[��H��dG�iO#��ى3���ܑL�r%���*�jZ#��'��	��6bt
eDL��㞒�-���J�Y�_4����0����i\v�՚-j��gɏ���(�(@㒿"p`/��r���rb����?sY�V�*-2`	����Z@.�J��Qz�T��ĵc�S7a	���l����0�����Yxs
@e�P��~B�d��bk��r�5 ,��b�!��BU�`KB�����|��RK�|E*��>im0A���y,��} 9f1�R�g��N�lt1���sP������,Ͷ5��2u��^�
��5?j�(U@��ﶲ�������bg�l�J�	;0T�.�%�Tm30;���7��1�����(�w�� V��r\��R�mz�=�#�Ϥ�����5�!�V��e�%���[^!S�W���Vu+i����T��#uۃ'�A&Tz��v-@y��45�z]P����8`�i��W=�,�Yh�XE���h)�g:X~� ��Tc��R�����{��NԆu�M�S�~op�A��O*t���>�����G�?��>Z?{�HJoYi��܅a>�L�;��8����Q�U��5��>aZ���Y1�>�ץȤ>�=ו���r����!�d�!�T�E�'@ZC��:	}[TO)wkh�S��\fl�.^�!4���A���,)P���PR�N�ۼ|�w}��0i���:|��2 �Y�O�*@�bTt$��[��~9�x���_�#��_�yn������[G+~%v|եH������~R�c+�-4��Z��/�i)k�ui��*�cp�ˍ�9Z���?�}�����e�r�:g�I�f�-{��D��+_Ũv^��zU���<���2˫��YB%�n�[�1g�I����HM��_����';1��?��9~;���=�0�F�(�5zM*��N-�Մ7�:���⡀a �?ⰋF�ٚ7h��w�����5_bV���B��؄q"��a��j����R>`�G�O��la:��#�������
,Cҁ8sn�PAP�c��7��y�#��y]=d���+���ᓨ'�s�O5n �<B5�k���U���u,�Q�e��  }�-ڲ}���v@��Z.�8����}��zz0
w���-p"��~����j�T}\h�=j&���M�Ɍ�<!}�u��a���I�pޖQ�о�rr�:�We�M�qjI��y����m�:�7�σ:O��M0����.��έpr��?��x�\Xږ�V'�	H��ELZ'�hj0!q���8=��$�������6i�(=Wrz�`p����<��K-��S���W�{R M�7�'��!��"�ECfk�����+��^��Ͼ� (��i�zn���Ȣ�S3���M �@#����m�Z�U	�C��G3 QӺ����l~Қ�e5��&'G~I�x�e�VD��NmC�����)8yׁ}N,o~QVƊ4��_�h������&�����)x�>�I�r�iV�`7ۇ6E{R��F<4R��c����IЦ� "��4��ɲh&�s���Z�ϯ�Jz~�������w�����,��W̾f�fV��r�,R��b����Q��=F�%.� *V�#�$����KK���o�r[�ŷC�2��N/m��;f��V3o���k~�ޟ�-�S�xffP�ϮG�r�C�N?��~g��;�"y�MLk��J�r��0��x��1T���/&���r���>�Mn�/)]�A��)7}E�G��r���������gN u����|-�r��®�m7�uw=���.�mG"�)�������ӴK9 ��tHf�B�%��I_���,��p���;2����l�T�u&X(-���X�*�u�����s�xdKQW�YK�o����B�5��(����
�Kz�a�3�Ξ��c)\G�ԢͼgXP��|��h(	�����F���ɇp��Q�h�<�|cY��y���7��q�������{+H�D��`dV"=<p�`kc���M�%���7M����zn�8K�F�ed5�$/3I	�[�uI�ii��
����T��h��,�DK�D��M���h�#{!��5~](|��A�[JU�y��#�A�
���h�ACR,��a�&v��Q��}ۗ}�U�
xq��t��<PM�n�Y˔�J$�p8�/o'E|��d��vS��5x��v_4����4��zX{{V)�z��P0��Ǉ��S��M�Z��JCc���e����no� �t�籍̉@�?u�y��P���py���9�����ե<�g ('�H�-������p�U#-�μ29c�4Q�3?:�.?ϋg�w��3n�A��`7\�|��4V� _��H��R��dE�#�K�/,/rګ�pȋܡʿ�!��c�B0ޕ���	�<I�u���M-���*ul�)��V�
�\��-��x��(���d� �-'�V�L��-����'�S�h7���CW��	�B�y�у�d��cԊ�ba�vp��İ�i�3�<e� V�o��پ�y:~,·��7�&�{�I���uK[�rw��u��I�1]T�&/��o�v"�L��Z��HkR���B�B�"�#@8�W8��`1t�6>(�d\	��meo���p~���Gw���6^��Xs?�?��D[s^LQJX�������Nf;q1�E9}O5\2м縃o��x�)��|k��lc9pS{�mS7?�T^MP�9�HB��v�/����_Z�u�P���5',�Ӻ��H�j$� ��e&̯�c%o{뙁�.<@B��l�ׯA��U��z���3�`OU����"�� `d��ijO�w�?;t2�:*s���7����bΤ{�ęl�gau��,ԥ��̲���2�J"���Xf4:�-����y0�ֲ�>3��7g ~V���lp�Lx|;�
��S�ŝߺ�Eo��V+�.3�2�$�&a�I�@+y^d閯�~\�а����c��P���ʻ�*�vE����L����Y��:O��1��H�������X��:"��� <j�D��8s�e������t��&��h2:3}�3�����Y���q�ܲ���V4P�����[@-�b���?�#�<��]yy)�_�Y@��#���Y7U�ä�K��Y�CnZ�/h� ?Q"��d�T�ꦤ�w�U�!�D0���6��� 	K�C{�����ti&�������62O$��Lf�M�>�j"�l�@�>�c�Fm��&�^k|dw ��ҥ |�P�b������0KE'�*FV��yPHL�w��Mؾ��\F�D�����5��P�߆8�Cņ��u�ކI|9:�[�"���x*�ԅ\W�,�꘎�y��P<���[�u����A�����)&�%���P�E�y�ˡ�g���z�SA���3�Qu��0�Wy���Da���lh���g���Z�zɱ=��4>rt���V��鶬x\_�s2��ɫ�O��Ԙ��n0p��O�_B�<�!J�a��xRU�=�˵Z�����?sf�ث�*ƿ�ɵ*�Q����W�#��i�y֒ *.�p�?��\�����ޓ�q���5zE<}�y�hg\Rq!~_)�a9��%`�#��ʆ�͓�X���	�S`:��2Q:P?�uV�R��`��V	[�l!_(:G%�ތ��Ip[ĆaBF�A|�z\����xXi�1i�J�����V(�8(�b��ź���S�,¦�~D�݀{����_9��1^��HJ�EZ^��8�]d�|�*K�`E;u:5(��4�z�Ϻ$�����?�X��H�A��9���{ Y&{�GZ�Ϲ#2��;��s5���-L�m��B���:2~%��tD����uU��O�B�a��=����EZ��|f�>�<.�������C{�E4��܁�؂р;n�/}`&S��CgAa�((U���o4�v�L�>8�.FxĹnt�H��>3{��<��ǋ,������9����#LQ���
��`[In7��ㅆţ!c 5��+r�t6ۓ����;��(�<:��T�kxj��y�}��ѷ�:~��YCΨ{���R�	�H��!�<�RQ]����<�cnX�
B@t
�z���;�:ͥ`ѝ�@%\T�i���ڈ�Ŗ����M$�I�H_�ǴC���3��m�Z�k�o���&4�a��6�}3h����6���J?�n#Q�����:�r��9ׂ^�$�Q�ǡO�P";��c>�a\���4M�a�-YAT���d~R2@\!�#@��[
��6���(	�=�1}t�@��=�?p��~B_z]S!X!l��J�E� ���Z�$��c�kZt� 3�"��F�O���,0��Ŕ�;��Ɂ\�u�{S�"��PΉ`��/Q5-���Cm�~g�I�K�S�P���Q�\(呷����J�/< ��R#c���en�]�����;�؁X�N~�S�߾n�CGf1ӹ�oR!�Ն/Pf�%�}G6�P�
��o�Lw.��ij;~-H6�Zikg��w~TZ<<)YY�9�z����#���<_H�Bz�]���μ��t��9���r�A�!��g�d+hUѿX�\T�Eb�b��!����g�_t���;��.BLG�FǑ�\�xx�o��9����)C�:~��%��շ��\a�(����R7\���"O��l�gG��0����0E[E���w��|C�K�J����Nuu�w4Z��,bx+S_P�(�6�<!���-�>cJ�ԕ��Z
@�������9F�j% H� �uȀz᭑��@��ԛ�A�3�P�m��T=	|�ۍHN՜����g� �*�<����X������^��h�Y�T�u�P5�$�[$0���<��?�I�ױ���B�i�s�մ,n^����i-�T�c�pAYG(�\'-��7�n���!��!]�{���?#�ԫ��P�ޣ�[YS�?�m��k.$����M�OAC'J����"�n&���%$�.��~��x�Y���96�,]ix��߼��a;&��	������aK�����ߢ%H�'�!@��M�||��7��8}�w�u�����6��%~�Wϖ�O
Y�/I�[�������S/��)�CL�ra�R����&���`��О�����0�ז9�_,0L�y�@�X߆.;9Q�Qvq����&S�֯�qM-X���:ɀ�%Q��?���	�@`j¥���Q����X��U�[���������L�h����s�M���/�sץ����'�+�0�4N ����BB�������BV^����8M��.)��	~bi>�t^,���{W���w��3��Vk�5,v����*��m��U؟��!X&�٦�\qR�Р�>k �lmk�{(qj�UQ��0�����gg�����2�o- R@�}^y���'G��`e��	��:�=�~p�Ҹ�O�|e�wI�n��c��=!R���	��2�F坞*L)n��w��(�p��l��i2��ֿ���_jG@���/	�g����՘�mνg��@�l	I|��_��@�dE4�c��i"����U^ӎ�\��5r<E�f�j
��x���Wܜ��ܬ_�|U��rNXu.�h��Ȁo�ܝ�QB�?�' �tA,r�}~�@����Ɣ�Em�s�/�Ǭ|(2(��?�TQ��5��1M��E�،M�a��ox��ո��A��e��I$�N��~�d�[�{E1Y�ʶ�����@f������T�x,�	�[��/�
+Z�;k�	\�Wֶ�NRw�Fºt��ͽ巫���ZR�kPK8ӡ-Aw�GQ�//W���RT��,�낡E�R��
L����s�'�8/k�Hpr�gUc�@_�eV�+�x7��I�2�0E����]I"�g����{0Gg�S������t��)!���3�D����`=ވ�>���g�}�̩�L���������Po,���t��Y�@wfMg��Q��؇0ʯ��\X�F��a������QD��Q����^쀫p��jPB6���#�U��D�����������҇rl��ͧ(����{�����=�_�uT�Q蘫�<O�֣=��P������Y��hj�6u/W)n�a��.X�a[-�2�>���PR���q�C�Ɣ9Z<�qHՑx#@�?zȺӹj�V(ޗ2���@�«��F��a�tطA���Q�x�W����H�.aD����c�єf��KC)$��An/)71U䨩���9��
V$m��������buwnzzX�0�-g�,���,tl�T̆����}$9رJ�]x�`eK+�,T�����@p#r�;=���Y>'�ѻ̧WF���2;�V}:�A&C���F��Q��78���8���8��	�<��V���4W�Wvg��VmD��@8{���m��Ӑ�c�p��=
��r>�e�:*Q�s���[������>��!��d���Z�y�����l*�H��F�`��s�['^�y�ؒd-��`Y�o���!��^$9���则�N�$SK�б��d�	g���W_�
յL��bt�>ч~�$.-W�jp���E����b����Lko2�ox|g_����g�-�s".����ƽ�_K�ǭA��:�,��Bt�)	���SSC��qY.Y���� WYɝ�w�]'��辍/�t$Ǵ�?�t<	�b�(���ٶ�{�]I����n%�t�-�gJ��J�kĸ��k]̬�̸�ow^P�^i[7�bdc`�8&b/�b�����ε���Oj�$R�lZB�-f��T�d.ټY'}M��җ.�[*e�V�ug�Uo��16W��$�,���M/LED�m 1*�d�_��?�"���Z����SL-�E�vz���y�q��u���zz����!�"7�3�������T�GHy���#r�X�	�Bw�Ndד��P���H���7��[���c�|�b	��>����Wb-���r�6gd��s�錖�Ħx>��=�>��v�9��C1�?2�K���
�ɵC16��dlf[un@����Yؠ4<v5��*tw�(O�3n-�f������|�+0�]H�=��Os!��e��_�����wL�6P�����;=Ϧ�)Hf� (C�������� v���,M��l��BP�����{�
8Ѓ"���m(?�rn=� ^Eg�n3jjzm��V�}�?�Ԟ������!�����;��I�X��0O4W��@h�L���F���BT���(��	��F0VNR����P��������y�O豈�2t�X�z��<���G�"�L�L��CL�@�Z5��)���;>��&9o�;ڴ�U+���V��T
�M�r ��|����7����{{t��1�(O��[4%l���!X��@EyǓf�H�Z�l���E�#L��_������;�#f� �6=�g�iЍ;���vV���(�Cw�}W�`S�A>n,�,�②!!��Xt�e?g�uq��>���C3�a�b��6^��b����ΓY�w��8��;[�UU�&(4{C�H�Ss�m��y�6�����6-G2`�u3�B������_��9�֘�����
g_6JZ���)R7���^��ݣH��n=�)9��|t�1It bE����,C|�%:���᪪T���[)���-ȉs�E�\�!���ܕ��!Z�M���S؀SW�>I��D�-�}r���Wɝ菓ʱ@��z�W��� �p�&n�qaj��5}"�ZմY�B����
\7�y��Uv��H�O�hp�н�*�}�(�J����_�(/�l�S���9�dj���An������P���/,�P*�^59yM?Gj2��^��&.u�I�� �`��3�_���0i������t*N(�.��V�^����g�;o�<@x)����Ą�)�`!HĐl���ܞ�������Ow���z��D'�GwK�ۈ��dڌ�a���v���ik��}cc/"!v����%)fP���E�0�ɻ3���.?Z�t��'lL��;��_2�uqa��JOʘ���r���������l����%k����J@�C��إs�*`�J�c6��
�넔�a��1$�ue9��h>Lw`�>=8�������nW��-M�f:��(�O���T)��'g�������̕0hh�T�)v/��x���E,�m�2"	Q;�`�6��8�a�V>���9�ͺ.[�xG�C�p���^ǞW��Yؓ�Mm,�)�I?��+�*���/L��������q7�)�Ə1r���9k��?�8����[{7�D���C�]zt3�np�me��	, �D����E�[��`��5͈T8�B����w}����<�*{��{��M��
:,�{Ȇ�X� F��#�����A� �����pl
"Uܦ�0�]��W97D��|/9z!o�\����!!eD��,�d�+�$'�H�T�[v��V�%�l�bh}��n��N뎩~�Zb���U��[H5Wb�l�T;��3������~�L��\װU�EcP����L2�;)�!�O�2>0��z�q��T��1�Y�/.��t�u�3!q� �z�7�?Q�,!J_��ga��x���[f�Mp0�:�VΎui��L@J)s��|](�+O��Lk�x�v��+�*"zI��f�=��~�k9
a�W�������!�g3��3&<���p8%l*�K���7�D��#' ��+x��ɦ�b�q	���h<�+��C}T$�$>���y��������e�1�*\}�yQ?i��a�+ȫQ�UR,s�n
�6�c�;m�`�άy�QN����%�<���h�̉Hren�YTy(�7�3\�N7[�%�#����J�co�4y�䯦C�C\�@��	�7�pt�n�b�X��usZ��+���ߍc"�mQ�LU>�I��a2(l:�x�j���&:B��j%)��s��ACe6�>U�z'���<��&�	��q�3F�р!�W��r�D7�]@��az�Z����z?�fC�ܩ�2��p���.�������LA�/����?~�ɣ��XXx�$ʪ���c�Cem��F��(�N��#����p�:���3y�#�����ɠ
�ӻ(ê�������~�%��g������EK�A�=G#�U�h	�?�F����t�6*nMp�[�-�x-����8�ꂲƪB���0��]�R9ă���f�	�*n2�ץ��vD-��*lږ���2��T˅��H��r���F?h�e�<r���@�Œ��)�UN��Z9��ܪq�6/i�S�����k���b�;
J�	D+q�����Z%�P37�)��=�Ycvw���� �5ہ��b�/��싺���wU��l�\�n�@37���I���}TW� ����2�(���?��h���p͜�='�_����P��$i�p���۾P�X�?�8F(�����XA���2T���@H�wɢD��OG^j��s7k@sp�+����i�����p�-�]��=|�L�9�a��xP:J����@���F�;���%Z���K���1����g�Q3!�UbqU�R0�Yͦ~k(b
��b����j��y�w0tJ�A��C����\j��k뉻w������Z�մ.��	،���邵�D;��g��p:3o&�,�z��:g����6$�w��9��?�S��9��,�K�\�5�$��ûZ�VUC��o^�ZЍL���$���
���FgnR'/����_ȂW�����hO�[u���,���~:��A���,��Jy�����xDI2q��N���$��)�+>�w� k
�#�L�@��~����n9ۛ7���[h�R���=fr�r��߾���Hh�gx��!�����~�w��H2��G�y=�)�,7�����+�ZdS�`�0�ճ|ԛ����/AN��,�-*o;�:�����1k�3*�QZ�9��e#.Z�U@B$T�Z���} ����7ԅs&�G'd� H�p7~���T��Kx�U��e��+�~_|@�F���]ZX�TL����5qD���Q]�Ws�Rb(a��.\�:�_�	���!^Ǿ��ȧ�����֐��&[�(���E��x��؁��7ߑ�ݺ�GUϯo.�Q�� Et����W�O��E��sË+3 �J�9,3��F˪dm�n�G�-U��i3��C�A���.���w�[7� �`,�[���a��r��P��T�w�,n��@cS�t�I�.���,Ց��t���N�+6��M�t��Iξ���54���w@�} fT+�����ޢ��0�${(�|͙�W urJ�`Sc���o���h?�㧔ǜd��%���kU�����h�eL�����6�LGU�2�w�G�Ů@~%�ïo�0��畮��@��B�WlԷ$m@I��>�ܒ�����T�rX\�Ua�#�L�;xv3@2d��T��ro�!Z(Z�~�p j��ǖ�
2�����T񳳙�>�I ؿ�C�7:%��	�i"�@t�ķo6�A/�,���  �Yl-4\&�R��i�l����W�P��ͦ�ї��$�^6�1��{�b���ϊ�8��8ȅ�c�1v�?�Y�Q���/J!���B�ks�X�#��Z�f\]���z�c�}����=B�FM�V,a�-UK/g4�b�Q��0��ŅX�T��4����9vS-��Q��>�(�3�H�sƺ��}a��3�)"�������6�(�^��?P^� {h����k�}�@4nHin��ה��Y�'NQ�HW�]2�kVL�R��[�q��#�2$�h1Z1��N�EU��@Th�Qw��[�Z?ыl6�A���A���c`��G3��Oi����g�:{v�.e]}��~Z�d�-5�n\��O+�T�X�0�D}�6�r<#����ct����F�C�V�r*ZDH%hM�Ñb4PE�-�lE��ճ�
�'�.$�<����/��w�A��dX�gtvN�N;c`���J.��R����Ǔ�_�L�3N��.x�:Ƞ����.Z�Pch��딈�7�|��Z�?�Â�:����Du~�x;�-�O����4m��<]7aol�tAo	��!P>^�[R4�qV��&������8�3(�5�j�)���ѤRI�����[WX)�LSKN��Uz �G�nd�PS��M��vԒ�c��E��X�|N��0�*���Q���Y��u!�-8!�N�����l�sR�;�,�����C����Ϯ���]	-���ee���:�咏�Ejc5Ty�a]i������I݀5��?�l�E�|UXDө�B05�����2��r69����ܞ�	�0K�D�-wsb#P�Y=E�kl�}i�ʣ��}r�;�Љ����Lk6Y*��M�k�k��X8�k�AH��8j=-����'s���O���.4���8�0%�jأ�Cz��"}6]��'��Bc5	�`A�^P��\�;�(a�{�j:���������W^
lԬ.XS�΃�n��<���\w����q�~��ߙ~(U���6�<+8�+I��!9d�xB&���!]�q ��o)�nF�(��&lj/�6�#��C��o��R�<��|;�.�qe
���Ѯ�CZI�/A���1&\iG���C�u�}>=�M�;z�Wn��|��7m�!�ՑS���'q�Ս��$\&��@6R"��#����s(f3����qA�s���2�H��4�7��2iN�F��[B��A��������Q��`�I�?�J���4'(�u�S��������w��D����h?����,�	�a��[�b�+�i$B�C�W8��^�����.�U|�5��P(��D���U�����`T��Z�	_KP9P_6ؾd1fs�Iwd���[(�隷��ڐ��U}�1�Xv�ɗ��z41q��Ïi���$W(&��k�~e_�#��FJJJJ��ͷ��od�`�Y�-XN.��C��5d3aud����ۏ��l�k��3d�|.��D�=	���c4�P-6y�kxhF��:b�ǟh�?��TJF��I-�u��?6�
�qX����:n"����x���?��I��R�ya�6@�c��s7�gYX)X�0_���J�f�cB�>��t�I�Q����/Q��%ϣSs��#M��k�S��J5�N�Jp�b���c$N����q�j���"|��J�K̩6���ej\�َ����ܹ*;�SEX���Y@�{���3��
v/z�cU"���g������v�?�m��x$*�_�V���=���6U��Ų��0�_?hG���Q���D\Jv�O��N�LG$� k�4�{���i�4 uD���T&�DC�D�~��~�U�`�"蔃O#}�n	<"7A<T�QnPע����^��G�-��.T�@ f�£j��?�,�޷2d���,�C�S�5����9��
� ��`�m������- ��g��m*|X�Nz���
uu�6�Y�V����A�q��J_���N�v�q#����Ƚq��yم<w��r
#dgCRW��fGy�	s�.`��,Y��N%�۶"�Hx�Z�4��G�$��^�(�>dR�tw�9��� v_a������S[,�&�j�d�4�R`����|���m�cr���?55��ր��3o�%D�ڌۜ�Hv� =��8/�]S
��y��>l/X_7�\�����Q_?�H9Q�xL ��W������|�o���5�����Ɣ��{�J"��n�?-]�Q�e��GgM)���D[?��:X� ��Y1�?c��%�b�r?|�,P�� �h������^)���� ,�z[�d��Y�j�h�Gʺ�繨վ�;�b��.���8�j3�\N���j�pT�-OѾ�t�I��A)��w�I9L��������<�'s�'����$���4Z�C糘F����a���{�e`��Vܱ�7LLI�L+]�I-�t�q�m),���9%��fO�\�x�Hࣆ�����x\g,��L��u�Y��D�,�<K��
�R��Ծ�5����T=ip6X�@j�t5Fx�q;�זK9r-:�~m�S}�P�]^��q8��ܣ��I�݈Qj9���_z�~�ђ��Y�祆�o�1�4��W��A��qC�����5�H��C#� XL�[��М4��%f���y~�����"F����O,���q��SW� (��TP͸�).�oJaEI�Fqbxŏ>� �IS�~ꐄ����f��]��FxE�l7�V Z ����h��MF�Ԅ���.���Z���'z�)I\%�n�ں�E���_���+<J.�D=R��m�[I!�	K2��ཕ������l��T
;O�Ht��/6��y�P����SV��6T��N� Ǝa��N&V��B��3ԺZ�H�O����~�>��@�&�Z0��Lb��l��.�����g�%����N;�J@�%XX�0���fN������b8��#��j�R�$s���> <̺�eFxY����<˰~jT�P���p�.���X���P�ǣX;�K���Z� ��
w�L�bW��e�� :� ���
���V�
�}k���N��h�m9�\��� �?K0����,yՉ}����>b-��4%G���qj���٭�D*�*g��>MΨ�]���t����q��N����� �^tl�@�����&<o��Q�Rx��k�`$׭�3��MDt���2S�y������&���[ �ͪcN�����,���Y#�D垖��.�?X:Ʊv�r!s���@_@	r/�k�I�B�D��x��`�����i���Pӟ�̞|���1��/��*��c6��ѶJ}����wd����6���r�&�5�rO��8g�Y�����,�h��X�a?;<��Y>���
P�ی^Ѷ�r�h�ѓ���bJ.�D�7A�3�����W"��_F���y�| j:)��������8\�R�r�6 RS��dV[�dI��|��OU��AHwZ%���|2�~Kr
.�[��3��씣�������_qN�@�̮i�q�yk� �<-tʩ+��5k��e��UY�m��H���/d��imL�7���t3U����i�Y�3^#ń��ۈ�l����`�"_ۨ�N��zr�[�j%�.zkRc�b=�y�?==��>,�i��{Cף���NΗ�ep��_*�Xd�3軪{.�{(���+|.��'3�e)���Wc�;!�9�1V'��(����H������Y��P8����r[r)?�G'�������ᛝ����@	�L���i9#1D��������܋�b�xs��0���q����i��uP�S���N7
x�Q��;U��ZɅt����v���l8Tx��uR�M�$nT��Eu| �H��o��{���'/�3�\-pF�ʯ�Y�m���=j��Y�`Ek�o�/��#���GY�:���SJ7]�O��|�H׽���pu�Y� �m��+q�K��0ȡQ�	�Fa�e/3��Qy���b����n�g�M�뺂��=��ũ�R�Imk��H��YhD�8��|�����p,#,x���_7����m��I'	x$� �����e�^���	4����W�:�!�ȣ G?��/%��3QɃ��5Cp��hM�e��ܤ�Ԩ�#N�J�{��ط_���`�Y�*��s#�Z�l�ѿ �0�3��Jv�C����
�e'��oD��2T�)@�/b\�D���V~9��������<��:�
�'_�K���BjY��4+�-������-�����y	c�KXo@nQ�tv$�q�쌸�`�(ڊi��3�*��d\-��WN�ڛ��CF�L��z����kd�.b����\|X���V�F���0^�-�f��2�$M��3M��m�@�hS�<ĕ��$]BV��^"�J%I�( %H�C{oՑeІ�3	i��w��i�`	7y�z/�1��+;���:�s*�k'����ik�c���Փ�*��L�ɣ�&��p��l��g����Qep
��%��_+'峈D���7_���ksvRǂ.�H󳾗%%������ĉ�MX��k�1C�'�$�y��-l]Ř�dcs����Gn�������m�>(�Կ��ʏ|�F,���-�pͻ�Z�D��g.����):�(�.M-Mr6e��6�����Hy���$��U�XV����g�.G�/	"���Y��1��h�;��0[F��20	MO쯜Ѽ���k�Ҵ:Ik�Y���]Z
A�P��X��ۚݕG�%�Y����<kB� m�`ғF�i ��b��7*��y�];!���,�1�|�^h��Na��K܄	��Jb���[�QH��I5�3�9���iS$��n��y�>-��;��jʇ�&��b*��q�`%�	���Is�%w5���Uf4���?a{h�4�@ĢL�N0@��ߑ��֡��Ė51ǎJ����*��d���]�i%�]U���Si���Ҏ����c���l������X[:%S����^0��,?u;8�vS��8	`�J��(b&���3�bP�&3��t������T�w��l-�1��		X����1���VZ�_
!���o���T��Gw�%f�R%P�èe:pp�5�x�λ�/f;LW�C@���uN9��v������;p�#W��|p+-�~�a'�8O�f�)�״KE~�����_�oV3K息bR쒏ۦ(m�*�a=�p���ԗr� ��o�0u]�T��j-��_�5�g<���y�����(�Ҙ�P.���7�r{��i%�k���9���	����A$�Y� ��- :�&Km��Qg:%�35锿I�$rFj'�>�]����J�,�������0�BH��0<i�N�>���U��lRȩ�!������h�N�2mzJV��ѯ�3���_��Y�8�N�/�4V����^�a��a��S [n-C�F�/Η��F;�gkl�����`BtK�c����3)���$WY��~���m;�t�3��:Ȳ����ix�u��� m",ZU���l���c;��q�e=��o>��Y�0hC�yo�0L7f��������H�6��
��"�E*{
���jl�ac��$���% ��pսW�����w���|6ѝ�r���l��s??q$�?tY,m;�S��~5�������f�UC�h�]�����>EoƤ>zT�"���1���g����R�r�#w��rJ��V3�q��sq�˫Mւ�e�rZs+R�Ġ��iL�fS�k'Y���ь�	�}Ҝ��s�}�k:\h	��r�-�-�g��@��.�*E����Dgݖ9�p�"4��ސe���eU��~����K��+=�����@b^��c�����	%�D[��Q�Gj��Z��v���f�rf��H�>�N_���_���(:��yy&��J
��H^8��j��M��LCF�������%F�4�ePJ����hW ��C�pS�c�9��	^�ׄ�P��:�*��M�&i��?��qm����`�sA�/�.I�l�x�k�\�:9J=����T�b�TI�HnJ�K�[�ܒ��G�g̠��饀���ߡJ?\_�ݣV���fY	�|ٶ� �G�����=z�u��=�R���S@u;ΐ��	4�J���Ɣ-%���Ϸ��u�:q�1��0$M��X�s��Ё[K�я�vq��i����z�r-���bP�<$���.G����oöT�RL!�7�6oZȅ��N�ć�#�R�W��j������k�H���m�����Jq6B�@N��K���I`�π�U�I@I�"��\�=�d�.��� d�h�U�R����G���#s4������F�,��#��s �Aı$W�,:AC�OLY��{�^�n&����%V��Hd� lK�7!l�?"�g�WQ�|S�l�`�x��o��񑍟��DZk�]��L���o���[�8�QoT���P��������T��z�맵%^<s����Q��8��3	�]���\%��h�����+|!l��T![�����M����u��T�HH��j�#�c�	殔�W�J׿,Df�q%~Q��x7���!�w�f�����,��ɻPA�H.�Y!��J���ǿS��6E���A�*��U�~��;y۴��+�Y0��1�`S���Ե+2��D�ˉ]�C7�^֞��C�KM��^�k�S�YX���\'C�퍢���V�,��"׽�
QzQ>����;�}3C��������|$��m�*hf>k׀�b�2��I�a�XJˌ�"(�p�u��{(��W]�Y`-t�n����-7�+J%Įw$,�Q�.m1=	{��5��%<���X�;?ݫ�kr�i���>����{��{�Y�������_G>��q��7x�S^3�^y��F)ω���
��'���0ŝ��,2��B�����Vei���ߦ��X�0�Rբ"��ı�4d�wv���:S�5��<�%���$���:����g���L�^3�S\<�)��V�P��0v�9#GD���AT����̈́��m/��mR&l�WP�]e
D�g/�*�l��u���&V��`L���������r��W��:3#����"(�p�y�MG�=�.0��}�o'dw�Wn�;��1�K�Z�P}�f*�ġ*� J��a�L7�4Gg~�J��/��)�m����GW�n\��AR���X�qp�d�����gtVq�\Z�a>a�ܤ�I��c��Ɍ�>J
Q\4��Y�el����l����Z5_~q��`K"c��km���*$:�n�1kT�W���u�@�P��^�.�K��ii,�@.�B�goi.rE�#�itNۼ�+�M_�/K'� U�KG���?`m�&�D��(s� ��ު�@�(BzB�t�:�w15�:?q���Y�z�蠦 �+Ӡ���9E��a0�7@�N���C��E��0^���$�P���ܸ�$�	��6�r�O��)�6����6Vqb��+��.?e�\[�Ɠ�"�]�����d4�f�zqI����D�K ���O�ҧ�C�Ԝ�Y��]~�OZ���K��C}%)5�	Ȼ�
��ޝM	 Gvj�W��t� �E�߹�<�Z�/(�$�|;��V�|��!XE��|�+�9��!Z��Sp�۾�qb��6�N�V��p��������]Q��-��r��Ǩ��3U�X�*j[��<J{}�e�aַ�����,{���Z�P��2�+F���
�S=�֝4��oC�[KC6�Wt��3�!g��l��A� ]HD�4��|���Wo*F2e�-L�%�^y�o��~�צ/�F���8)���q��B-�y�=�S�Zb^��A��3����OJe�O���N]4�F�T�&��q�+�v7E;uR:D��� �D���1�'�����sԻ[>�n�s|�p�.��@����"�������[�l��iB(��w_\f3�&w#��%V��/�n��k��Lb�G��	�~��~c�"a�4ӎ�L�PP�a$|�Al�,�/)J@ �	u�?*�8� �*�n�rSo���8ˠ��?�� ��8V����@�6�^z�g_x�S���s9/Ϯ�^RHהӿ�m_0��� 2a�O���w��ႏ31�;��U��	��k��aCS��H�J�>Ȭ��B���j2�jp�i���h��Y��K��5[�$>rgs�J#i�u�zy}�v٬�\���⌋�+��_p#	�R����O��z��E��)��e~���)��߈�e�������HcX�z����p�Qm�n|AM2�%�h-��)�g:hM�`�-D�E/�{�:�`� �e��b���'m\9�>�􀕙z.��S��	e{|�'�T���6aT���W���Q0�A���.���5Q��>���2�����M�V�	�f�a�[����A6�nK]�m~�0q0����8�ǜ>�T(<���#�V�4 ��Bd؟˼*��^ϖ4]5!K�3�� T�������g�����\ݪ�"~'�@vTOd�#O$�S�����$�6= Z��5Cu�$���C�t27WM�>��_1,�`!��:j�t��6�m������,��DN ���n����P�^��E���y�\���졄�k�%|s-��i[8*�!�>���x	C���Uv�G��8\�J�i�ʧ�U�xO)2������*eWQR�J [:�h��@��z����^\z`~�=�Ԟ�3;?+��s�OR:��5(�U֔��`���=�7{*�t��TՃ��R�!;y��k��_�l��`@Ô��H��/� /�>%{H���G�����0-�Δ�����r{���ԍ�4��e۴AB���T����m��QY��ˠ�k��2"�zH1��;�;�� ��x|J�X*��@��̹�	P-Y��a�Y�5���L�Ҥb���0W�Ѿ%8]�F�i4�cʮ�v�p�)R��}M�Fmo4�D�]���x�l����G�N��n�f����㍏p�o�� mF,�/&��$����Y��Ԃ
X�$l8piA燻�9����y1$�ǻ��>�!��~2T�}kA&�/���@�F�Q&�aFw�ԯ�:��_��a�3�a6����ru��.��E�M��h4��C�"Q{�:��g��mkdc	|�=�Ԙ9J�؁#�h]�d�~`��qY�	jK:�_��T���<+?o!_U_�R<z��	=r�E[𝓻ǤE�=�H2U�bq�7��5�'���|�-�1j<�fYpG��i�i�������%�L��W~��o�� �T��p"2ڇq�b��U8��6T�i��`�Ě�g�:�[�q��ī
�Nu��ڱ�k��=�Ry���7�������o�m�EICf �Xe�n�u���(�m�=��Uh�q�~�7���I�j����(m&1���J��2�Q���4�gc/FO�kFl�� 8��
��oLG�����z���YZ��Z�\V�Ea�|H�?������=�J��{�5Fq������`)I��`7���1e�q9�D@<v��BX��v"����������-�9��6]]�͇�ϑ�}���s��t�M���'�s�o��(���:����!�ǰP �7�ewW4QFb+��=#���Bn��c�ő������'��y�o�� �)4on"��I��2����
J�B2��m|c���ag2��r��\��ՄI���"�r޽�}���.�	~�_u�Ϭf����(�F��?�ל����I�?j���G�w��r��GN�f��P��� �b���73Շ�W{�Sǐč�v��1�.���hQ�z���J�/���x{��I���᫹`�Z"�h�y��ݴ
�E�*f�{�$h!j��+�`�:���݌.M԰���J�!򞀊�s���v!�>2� 9�t���[�W�z��(�,]%��D��,�ķ7��3H��^ ⭛�����R�5��"��|� ��wE1�2,���C�@T\���.�n>0��J�I�|�ʹ !��,K���`��!Ja�ȯ4`�繄bg�wB$��tX�4.=�t YU�����혨%�)y�&f����&~���VM���`�G�#dK7�6ܸ�6Gb�ɀ�ٶՈ�����
~�,=%QÐ��%*fkĨ>ȴ%�~���>~Dx@�=x�&�!���B�Lc����D�#�u�8�c��?Q��!��z��!K�(�/a&���l�1�nߧ�%(�{Q
���K�欄�`y=D(���:iz볃Mk�(W��+���6^O�K<y�,d�-��)���Ӥ$d�˝dP���M��]���pMK��G���_�a�iC爓���GĹ��\�J���<�nV}Ҟ���ow �;�PF��DA~,�T�粳>�K�AJՅ*>�t�k���D�1;��v�d���&�-���>����EO?�CP�	�w|�\�xZ҇/��Cr�G�	a�Q���_Brf�����b0�
����#��"u4\�Z�#�G�-��2{��qc'k�X�Ý��S�Y�8,+��h�r�sKxGv�E�͸�1-g����fD�a� Q<�w�O�mɦ�ŭ�r�=X�n�O��6�)����΢f�Wc��vEv_�V,P�$�d��I���2oA^�=V�A�o�!�@ɂ�+��X����s��=1���.R!V�yx[��wd�aa�i�+��Й���C>B�C��`uШ��0�d�jB?��:ί`Z9vn�< <��TB�����
<i��ҕ��C̫���Q`G:���"���A�Ǩ̍06��@�A��f�Mթp��p��*+��Wýk����RDa�x��۠H�)�]"�P�֎lJ�}ſ�M!u��+���3/hL�<�M�J�JW*�>rK�V���w5�8��2	��k#\�*�2r
]s����^|��|٬�R?)1%�gBV�(�Si������������o�k(TT��E��?}�KQ�z�==����c��+�F��.�U���ڊ�E��1P-����}FZ�d���:�!F5��س�+-t�N��H����LvU��ݱt�G�lǊ���)&��]]�E�.!^\@`�[=�u.�Fژ����L�E'��bŎ��`{�V�Q�=�G�w�6M�s��c�+苸�?g��jj���2_ա`v#��bMV�M�����Еi�����'Z$l�tT�]�4GD�G2�o�p�Y�.3נ'���l=����@��ډ��T�F�(D��}�ʂ]�^�On�-����`��Pvb���u�����t��]Q����ֲ���?6R]�hGq"�������>��:�l���qO����D���x��
��#
l��F��L[*�/�Q2g�?2cZ����_ ab1xe�h�%�,"�����%�P"��<�� ��b����"�Ye�3��0=�u�՜��(RߘZߋ�Ws�����,(�ՕI�$ӯ�/��3�$_P��mH��
�pVyUf�`jF`q���e]����Ū����ě�%�m�E�G��%:�2Q�v��u���U�hS� ��q�ax��?7q���&Z��s�Q��n��h#��}�1~��[=�8�Mj�(~h��]-h>�6�0)��W�����x��F�ܫ�r6·|�j�X���\9����8�(.y��J�]JL!�(���ٽD@%���YZ|+>����.mL��n=��O��h�e$2$�9I����VzӘ��%*�؟⡥�T����#�c�툅�<i�CT�Am�_����_��ʙj�CD�;�������d��04��bڇ��r��۟L� !vl��kt�:5��o1�tSէ��ɛ"#(d5E7�pfa�b�fv�/����v�S�k��0��i;*�,hs�	|J�k9�?��T�O��/�-�3G8�0O�T��_�iy���-+��f��4���0�X���*=����vts����*¼e]2̨��Yq�����:���yGC$�+�\{"�7%P `�5ۗd=^����Pn�Nc�|Z��a��bi������zg%�-���毴�W!/�c�4`���s�\�#�cvns����YU�*�ⅈ�Gmj1I�4�LK����e��E<���lA�0t+�wF���$~qr�i(�f_�U�Q��Ey��~~md?��o�|����0�O3ǋ�f\0�i��)J'�1N�V�7��+E�Db�?{��v�U�졺S���Xi=��s됀YH`֊q�!̝zgoì�q �u\%"�`��7�t_ir4Z{�"��b+��t�q'6���1B
|Pwgk���,�ʱ�E�	Į�ކ{ N��3"2'��_���a�_�7Õ��\�����1�ڥ7]���Z��4-�4�W4+�E�U�z]ţ����^�Q���k�4q�]��V�\�:��\�ҏ�[V��{��>w�0�QBm�)��	���Y�qk����'�7�蒡�/`j��S���lBS` ���3x�����H,�,+���cB��wmN���r�;u{HL��A��t�:�~N����y��u�fh��`d�S�DYx��+���:mܞ&���'��@i}�c�c�I��a&�5!wwLW�8t�B}gh@�o�������N̤|�jj�F}��'d�`�.����6��'ABv�O�d���J��)�
E�;�/A����<[i�D��C�댝R+�V�քl>3T��Kñ�)����H���ł:y���j��"�A,(c��%&��Y%9�{@����'�y���o�=᭕�s��t�a!j_=��	&�G�(/�D��4�O�`D9;6��"�t���4XH�7׋?hl����p�ֿw������������j"�9��jБ@���3�4��-����>J���p�+8���3P��7bP��K.A=:k �@Y��g������Kk� .�Z"��9=`c/z�Y�ǂ�V�*�<�	U��>��tTb5�×ƗĊ�
����O��e��D��q! �׈��G�F��'Z/"oC�z�f���Sl��	����D����s�1�����!R��8e�E/�l���~b��u�4���!M��b���bd��B7�<7���m��[]�:	��N��b�֊N�D��e���ߜm}B|4L��zj9+/�r�bD�<n�Q�Xl$�B@:McB��Ҭ��:���4�	�ǰׇ��6%+̅�V-�|4�
��5�@aKZ�C�gyt��P�C����;��|�jh�a���mW��1C�Y�	��^��1��f-uvjH�Q;UAf���wn�K���wxm�ĭ)�O�%j�����pr�C	ٸG*���T��7/V$�.��h�7�����2p�H��O�%A�l��+�u��y��,-���႓���X�� f��J	U���Si�'��q�4kj�"MW�����ށhs�+r�Eĥ�	��H0��1��@�:^4G���A��a�B+����Knx)Tt"NI��v�G�?��ZC!1������_s�aU��w�LS��Am�ؼG0���~N�[OO%��JR�WZ��c�u�
L��3d_��kXB+�x�FK�2�ⓧEs+�]
<E�U��Ĩj5G�6�\҆:&�:��=B,w+8�U� �5�	��Y��ӛg�J��Tu��]�jG�pC�Sߋ���X�,C3J<K��gj�K���2>��8��	�ӗ\�0��wuU��w訐Ae�R��k�D�x�}G$z�Ne�Uv��0�C��ˁ^d���kK�+�^�E��V�[��$c�N8�����
�� 8���i,K'�2�%萖<�2���@�`R���'FbꟆ�J��+�<�Q�hrQ�3:��Unm|�iI� ��Ө��Ӑ,��>���/�e>�iJLb�Eb)>���������, [�S۫L�	Vc�%��=K��ܫ�֍�T慨���[J<�$��%"ݝ9䩔ԆK�'�r�ϯ�Ԩ��eLH�hDz�E��Z�_�ks?�r�����Qv�����*��/�3��$��ް�[\����5|��|��?�>���� =��χmV,5l$�I�����1ϓ_��ã��xM��6tg�s?\�������-Co5}���i5���W�MO�\뇊k�@p7�g@��<����}>�,���b�ua��4b�$���l��A@��yM���+a�ZR��}@�j���J���.�J�b�Ԙ�ץ��ꔮV�H|XQ�9�����V���>r���W�D|";�'&-UT�"!���>�mv��
\��+l\?Y`O�Ȼ�G]_��"��0 �FH3��&6����c(49�	ꓰ������c��Qx���}|8Sd)����Ѹt�d8L���&BKXi�a���ɺw.Ok��OIZ3��ΘVy���2�B����ؕ?9�Tf�܋��|�B$>�b��D���2���nJ�J��]����5�/�Ï�����<� =jǑ4��yq]�0Ǯ��f˚Z�4����ے`'I�*3�T��!��ڒ�^ب���Z�a��>�l����o�A�0���n:�!���3a��Wq�1Aj!4����>�M������@��b�/����B!��8�#�kmM�eC�Q����?:;{�~����l���-�O����+XLv�ՊM&f���p~?��)�Z�Zc��72vH���m��A�&fp�CRi���nH��T�J;���2�u���
J�)�F��)��N+����x��v����[ Y��rv]���I(�Qj�XQ=gg����NI�*��d�SRi�$�����+� ��V��F�-u��a��B�k��O� �<�RޢXXoG��8ᓕ����UvW�9��S��x���ZN^j�G0g~�e��-ocG�,E5o��$>�KEo���W!�N����E_��G�+<���!����&����>it�%��,�<�4�p)%��|+SUWg�����8���Q@@N��ͅ� ��	m~#HQ��l�-���c��Z�,���,Q0G�Jc� �����-W���4�9�����ٙ���K6juZ�PI�<�S+��>H�m8PA�����ԨV����cW���j˷'�0�i~�l��6U���wuq8
���J_���G2Ψ���پ���C~R��!��Q���󠥦��ɚ�<[f�V(O0�M�x��n[�R3�"�#N���/!��Q���OV��;��A�p�-�O�b$���~����S�Ʌ�G�֐#]]0=�� ���kY�m��b���n�m��L����U��e�he�-�FoƼ�,S�(*� �T2Z���?IV����z,�wiE�BO�����n)�U�Z�#'σ�qO�I�c�ߑsd*Փ���
G�z�'}�'�
p�a5=!�����"O�N���!����u$�n"��[[D�T;�D4��h�Fs�ǅB���뀆�Ǐ��O (���@��VrQHox��d0����y��]��yvB!`�b����o��X=H���]l��V<���	43��y���66���vgY�rA�6I�?�R̖��+ :��P�t���+�i�$V"�&8��g
��\���2�)�de�Τ?Yں$���S)WQ
r:�)=s.��]����b��6كdb�u��J������`��7bhy�X��j�aX�І�kg�V`Ojz�������-����4�oM�K�l���wE�A��B���<�ބ�`��6dY	�u���=ڰ�g�RW{��2�9m��|����dY9=c75��*0|���b[)�\���W�U�E-���Zi���d���G����")�8�[& �^1�����C?�I����5���u�)ٮ�C�jS��B��:LA֦�L�W��g&����m�h��y�n���,<�?�0�'���Qib�T�f�@�B�����h��#�7+��+��}@Yq��Bo�����j��X��D�ż��4`e8��#@�i6�)�D^8F�R2�l:%Г�z���٨��lr�x7yn����P#��?����ܛ&���Lq�P�O9-��v��2��%�]e��PZ�7y�Qkk|� ��gNv3*u�#i>��	��o���T��7�PE	"�#|xh('��LT�ȀȚդG�v �O���b#t/gs]�X���"��g]tu!0ƻ$�� �Z��q�Ε�e]�(�& g�?/���෩o�PnG ��Az;�E��+�Q.��~8ɉ���lO� ��=E��o@ ��Ȑ��k��r��Lm���p1&�A����Yb�<�_#�N�iW�<����.4h�*�䭘�̏2�8���>d�4ڇˤ�t�/�5�4`[��,F�'�HI��fa�ڂz��vS�'5�%�C��*QPMI��[K�<bO�,֠j�K���u\�A!�W����,��#<�;Wҽ����#��R�FK��PVS�0N��jrO=��Wތ�E���P��q^Ԭ���B<�z�����d�s:X".[˷�Hͮ�.�e���s�������@�4� ]Wߑ�+|ξ���T��7��8$	��]��+�f�2s�s��IhQn���:hev4�N}E"�H �}�G�zY���U2�����Q�l����Z-��� ��9�0?vs�FEu�����_p��Li|H��B;w����bth�l�\<��
�َ.��t;A�`-�:-��lL����ŵ���G��9t�g��Z�<�m{%.t�J|�|&�gq _jդ�?M�}&��5��`y:/���n�pţW;;��Y��Q��Y�5��ou�R
��]�R~J���;oT<�H��9%9I�ָ3�ۼ1W=</<IS�[��k�������M3!�N��0��RuK��k����J���ɦ� ���4�N�$)�FF	a��b���i�q��[���A��"8�/[jڑm$K^�>r_
����(��"�J�C�I).`���H���P��^G��+�����bz<*�?�8[f��E�A֒r ١�`�M1*���/r
4�T�5Ӛ�Zѱw�䢵Y��tb'Se$�H�i�V^�x.���˸�1�x��#!/��L�u�C2`�!+��&�N��ZT<m�۸4+�8eKE���5���29uGb����#F��}+��4V�v�"͑��P^�> ����*y}�"�cAvf�]6�����Q��-B:%^z*�Z�KSt��dZ\s�Ez�2s�?��N���@��W[2�c�w3D��*7����^��O�oϤ���zΦ�H9��Ǧ4	�mn�֗W����9W�"�E����.
��6�3��g�5 ���e�?�I�;�L��L���ܲ�z$sq�CP���]{&����Z�-���_zb�ѩ�����ܯ�A��\���UX�n����<m�fՂD���1�F���
�׳X��E��s��G�*��~ۅ`��Ѩ�j��1.��;7��l����ㆇ;d�TT��.�;ý��S�TI.�,�ߠ�b����c�BG���cra�_�E\�h)*F���;`;�/8��S�'+W����^8��HOrJ#�a�z�Zy/f�e bw[}��������]����B�z":"Y����k-)�B����2���jN�/��@��ڜz`)��a���N�/�Y��
*�q��jfW'�s(�<c�%:�4�M=�D�B���7�_��؛��`�g��w�k��nłL���U�OW";됶�?��g�j�*:�]Y�a�����䞅�@����V0C��LYi9гn݊����ɚ�L�Q�;�0�qh���,EOL�b�T��lV��=�g�o3�Q�T@�!ɂP+�Ta�Q�I��[w$|%e��@���V�c�Eo���$}^�l����XE�S6n�=�}G�>��zfT�頰;N�B�'�	RaZG��w�_ i���L���������4E�>^IRҕ�+oO�Bt�k|-LHT������Ym:z��AT�Ӌգ��Mcc��[\׋sF���i*�G!k���}�uO��l��'����:/���c�m$U���m�ȼ;��E�D��lM��Y^���5js ܵ����9�5s�ߞS����[`y�$p�e���,#sHθ0��5�5O�eb
BC��־L�������e�b���#C����K7&@���^�	��1�+���~R®����.�(]�~��,�p���).��7��{Eߕ~ȳ�t���sڡ���%<G��}�3���j��fg�PR�K<�����N�)��UO��w�1�RZ@eFj�Ls*��N���N4A%et�H'�BNm/���qY�V�
\Ǿu�-EC�� _x@ݡ�.m��ؕ���@���iQ��S�q�ҥ.�t :��撂@_�b����!��`�`H���t	1�����>\'kXa�xB��~T	�c%��Ab�c��=5	ԏg��Yۆ�k
���G�q�&2a�Q1�I�p��3����wԁA���~�{�sj�~����=�=r��U	�gc͹=JVΖ^4�j�O,$� �3��~(��6��"0D�l��QΑV�Fo��_,ӻ�	�����?v;@�<����K�K�q'�z���C�G1�b�)��hn#`G�ŝ[�I�I�p�����`� �~OC�@2rw���{=8��EތQίD�S����v��E���n�U -�<%p���k#ʽ��K��(^"��HK�N����U�R�$��Qߖģ6��C#�%%���~��E ɝ�$�rtc;%�IV2�)�1�����0T��rt��dHh��@(�!��0@��4���,paƾ?quh�YIA^��*2������rB���B۸ ���Ԉ�K3�-VV?��R�q�Nnr�,Fb���v{����x�d1��@��-����aza�M���\�9V�K�t�D.�1�M�mq�0`�1��C�w��Us�hh_���JÙ�y�2��=���ʃ]�U�\��f��&!X���|9;��xv���H_�8t*1)L�Ĵ�ɿ���W��:�o��.$Nȁ�ԋ�Z���s��8�������He��<���C� ���R܂�QT���Z��\��� �b
UB|���B�s�Y�Y�lY����3�3X�(0���������Fg�vr��z�Y�7Z�HE�KI�z�1PqW��g�>�Va"\�S��iDŊV"HOf�\}X������(����Y9�cFc�\�:_���)�/�^_�q�(���?�(�w[�z�w=�Nz�D [��7e�L�vy������@�=�q�D� U�?ϒ���eL����fi%���JF71 �Z3�]՜���>���y}�=#>��!�o��S��`�9�� ��B}��+'4׎��r��.CA�H!�jgH��R*5��G��g��A�Һ�����4�m�������P"N������.�o�"��l7�ęi�pB�fFj%.T�I|:�����%#إ8�uwg��ԵoZ�$�~3޺�����ӊ�y��-IbI����+g�j�\��VC���6�^��w�~�*]@�/dk�GO�K(�z$J��1��J%oH"Zi��q��vX�vYA��Xaw�����U��y��i|gH���g����GTjϭjh=A6Hd٠]�[�մ�ˢ�;f�^1 ]`J��_A�a��]]ƢIT9=�⾄Suj�l]cMWn�?��9|,��l`�k���1�z-f[�%J�=�2^w�:�fpC_�#�E�HkHR���B8�`lZ�U��r:+��.\��EɀJ��FKH�_�e:��o����[�-��-��0Q�$����EoVP��!�J�>��.Z��Bua%Ԯ�`h�g�/qb��pK��[\O�*�sD��.�N�]w�7j9�Sc��ּTBu�擔̇�xOI9�+Tpc�X�;���n
��7 ���=ٿ�qnδ6�ѦJ��v�<6)#.�#�(�UʀR.�G�l�o��1�a@��L0����X���
�A���b��Aun��V�^�ʵ�����I��aS�E�Xp�b��Ejr�jj`�c�5G���OU���F2M�yX�pa�^���E�i}�!�?����IB�Ur��)eƀ\^C#��?#.�a�L�ջ�dK�̒�!p/� ?�y=��Hg�B[�H�y��f�*��~�g�k%�nɓ�T�w��2�9 �c�y�=�v�*\.��w��iD�pGL�f�rנ�t3B쮞}�E$�XLt�W��A[9��	x�,C}K[?�며���b@������{��~���lan��مA�bQ�:KW0Һ.��m���	��^�M���'i�f�7�k�3'�1�Xݥ]eX�&a��W��:p��VI^:��G{x�)���-��t����	=��c��j��}���U��O�p-i�\>˧x���*����s�i��y�x�����������A���N���NQ#e���SN���P��_A�{�ż���Ԣ��2g��/���{�0���lj����L���e�9F�F���y�E����"����<�6t{&���6��O�"�ק�I�ǡZ�g������&�����F���;`3��~�X"�p[j���E�#?m�Z=Oi����$��I�k�����<� ��f+��2V/#�
��p�9�#��r���G�Hq}]��?��½����عIx�td�{y���P�
:e�z`8�k�H��>Մ�[`���6uL�o��G5��0qL�B`���А�վL���NUR�����H�����4��D��1\!�c1�_Q|鶚O�8��?[�rt)4�c�Me�*���oaq#4���;8F���T�}N�y�J(>�A�+�,`�xt\��s���琷���Ђ�[N���h�'"���_zڧ�T���t���r��Y��a����	8�J$��5��6��?:1<l�e���-�t���F?��,�8�a�?���Q������>$�㷪A�q����lݮ��.�lI�V��YQ�ͷ�vO`�ڡ��(pR8o;6�L,�dX�!���G�Ô��w��/g���|��b��1}�ק-� Q+�!�!��K��n|�"�hzB�����͉WF��1N�f� �.�9ЦmA�
~�Mb��v��VR$�?��z�ǈ��cw�Ѯ͒�}�4Ca�l5A�9���x��0�#�I���L�D5���J��TpL�G���#����.%��=�B����df�$!� ��oɾ�{<ϠʯJ^I�(#T�s�y��8ŝ�tf:�Ø�ϊ��ɿ�(���*�o,*S��|9<USy����p�9���1aa�觅Wz�U������}7hW��V��=D<ź5c��}Wf�	�����Y���ɋ�(,�@���>�,���N��:/�OlqE�� ��`tn����`�	�o�π�'8��d篵�mJ��K��4V��g]�j�:pF&�'��=$w�Wn�\QƐZ�M���,���S�a�~�@��;��:_CX�TLρ�v+�k��\i�>/�ɡ�����J=�c���-�QV��20z]]f��?>O�Y�C��� ż��zi٨���f[����-���ۣ�p��]�kg��R=R���X�{_O����>;�/�_ǈ(V�a�t�`��������W���� ��9$��-x�f"-�ޜ��f���2�u�{�8�׹}�xtnJe��)S5(���`k���Ku�*�+rHD�?�Hǎeuz.Sfo.��50�8,��-
ԡ7|o6�5��硧0���Eas�4��E���
�
W4�N�a�R+E�Rc�3q������?T&O�{K���L�/�X�����	��E�l�Hr�^�@�;>i=���x;��{�H�
�࿻��A�L����pH1rA��1m_�.Y��(��/�M��h!�����y�iԚ�.n�۳	��V,�|Mt��e�ጋg��CB��O���R�d���m��6������Y�r	�5GR{a\�<���k����Oہ0Z��d
kԀ���ě��{B�O�N]�;TA���%j�Ob�M�0\��aGH=	�鶞#��XZ�XJD9�c��x�ܣd��������i���:<�!�S��v��떿%�YW(��������
,c)<��(O.��vWϏ�X����$�l?��_ղQxs�۶k�t;����mE�(R���m��
�:D	�2Ľd}��y�Ɏ�4��F�˥�1�TFa�^��*�@�|�~[�C8������h`/�M���P|>2�
���ӫ� ,�����4�VSz��
k�j��Kι�6)Dl�:��ɯ��m+���B�
����D�_~-~ҥ��	!d8�;�1GQ��r_k:5�}�~�;^�K�J%��C�#��=���W��ސ��Rꠕ���)�]�m��8�3���a9D��M���h����~N�N���Ӛ�_̳���	CG��X�~�{{S�%�O�nqC�9^<���Ѻ��>K�C�s-N�/�8�!�ҷ���a1\�oY��Z��w�Q����|=6&���3F,і0Dz�g�	�yw�z��m�}h�4M,��w ���AV�I?�h�>{y>���_�賧D&��\9��we�SL�"��Gb�n��3pQ�j�� ���ga��4)<~��Ɇ����[�:�Pw�M�����D� _ғ�8J�aKԍ{�F�ݭ0�aܚhW}�Ը����B�ǘy�))у*��1��7H���^�BvL~�z�pJ^d�+�3i�+�ҢR>Sp�z!늅
T�	�]�I��j�n��M���
T=�NP����q�k<Hȕq�x8��^�~}>Ԅ���S�Xe������c��XAO���L��Le�6�Y�@�n:?.&�Ib�UY�x�(s-B�(
�zRd�fLnI%p�%�Q���>�K��/8&�P'�����
��W&aT����_��4*��e��d7�x���.t}��_�zπ`�Mdd΍�_:v؅��Q��&6����Ӂ���h�_�7V��g�bЅrc����Q!2�}�*����2� �����+���,CawM�K	!�]���<�0]���g�y�QS|FC�d�՘+e�ʴt����a��ϼѿ�di���w.��;d�G�EP��=��W���~���YOC��P�}&<9᰸2=Fd(�a�6` 2@o�.�,�4�2�$���oy�_E�G-���"�Ջ� �K��`}���eM<�!�Co�83��s�zx�����f>��T��f��K�����G��P�lk��x�b�~C4�԰���A�W��D���g�m/�WYQ�O֯�����io�LF?DO�Z���1��@�<��C��]�+_����~90z�؎��]��B�},^�'�
bǷ�w"<���8����S)�`J�4M�+gB~,kwD�
�k�\;TG7���_h��m��5w��_�n�+$H���Q�ߖU���#�H�Y;��.{�������.��qw?�R�9UU�_aD�)�o<����-�zlf���\�ivc<�d��. �0���|x���$���A��P���A�>�p��U�W	�}ˈ�$�K�*��5�[�D4���S@�s~�Te�t��P��;.5���l8;�X��H�4�J�I׊Y�
 X�������.�ޞ���;�*�Y���������S,ra��Oc��r�.�����U��8�����z����,c����U%��	��ǐ6I��fH�rNH��~g~���+a/��^ _��Mk�p��-b2��B�������5/l�O�A8�ӸŃj)3�琯��M1�p����S��?8%��B�~�B�/�·gk�Y���<׀F�����/α���v��H�|A���ӧg���~�\�ZB�;���T��M�}N"[�&%�ɂY�G'�����c�sL���֙^�����q[�����s��- ��^c����a��B�XC��\֞�Z���B��&���D �A���N�[)q���b����!{��Ib���K'x�g�K�[��I|8lsC����\�utT5ꦅ��|��w���ϰ�!E2�[wh$�T}�D�9������ߕ�L��}mu�~�:�e{Q!ȧ:ڈ��
��,F��D>����K�9�\^����z�4�{k�9 � zBƶ�X.��mJ�5�����NJ�m�1݂	�4
[���;�[�؋�+�<�8KKs1����

��|���	�>�����u�Z���m��y)v��ӫ<���e�����4�B5�$��x�o��Y���{-,E��B�57��y�)�۝��+��4W����S� �]~�o�U�K(�K��+".�O�
�|��-�Zx�SS*�Ttǫ����L�M�AS��)�G����| [X���$�g*l;h�Ӛ����a�o��i��8�x?Lq�!	%��&-�
��Sj>�����3�l-a���d��7eӻ_37M�5���(
�j&s"a�bωC	"fG_ǳ��(m'��<�^�@ �D	>@��l�~�:j=���ɠ������a�>B�;�K�:�|�q�EC$a[O���yAY�SB`�#Z���(p{�S�L��AX�U��ޓ@�*�HN��1|�
�1]�m���/����Jh#��[ʌ-�_�,)ӍŦ4[����$��@�7��"�l��7�ڿRr/���c�D���4A�u��ż�N�����^#i��6�)�q�M�IF�DL���0��z����`��t�@	�&F`�X�m���ݓ�s�K-��	+�[���1h���ӥ�����f��!����V��oH3)��;�u��f{�|/�L� ��I��2�wlI�|(ŕ�B��U���	���E�N��>W3ɺ�'C  ��I~-����'<f]�k�Ω H�0rH8S
��� ���&'�P�i�t����'<ѳ��u9�lYx3�z��.�Y;,Ŵ�on�7�rt�4��R/B`�ig{�^$_�]5��@W[߳QI�ʛ.~��$��z8�F�8��qW��eSY
_m���}^ܢ[��+�D�,�f��d��_y��#���̎��Ene�����
�3�,��N �Zdv?*���ҽ3��� �z`Ū��6���w�un��S�#�bmC��D�w�|����g�&Ss���T�z �s` ��I��3����;�(/����wƔS/v�6�5]BR�yʲ�D�Sa�*Q'�Gq��׊-a�������/�,P���5��gG'�0J-pl���%��M"��e3{eQ��Y|��ռp=o3�Ez0�~���$}��^� �/M6?/����k���
���	�;��7<�vC4;�'�m��Vɗq=�r�_��3�Q\��:a�Ҁ�~<qX� ��Nז��YdT�s�F���%}<���A�{�ݩ�x2��w��Ǧg�*qu2�π�ܽ��uMy�By���p��<�jF��O�?�+>t�B�8D�����ޓ���{D*�V�:s��-��/L�ȏM]������͟�Y�@2�O� �AZ�%�h8���%Tk K�����`]�y�]\��2���trlPHnY�@s!=��O�+�*'�j�O����%'�N���|��0��(��0Z�_$�|���\D~#f[ �w�(�F���H��Җ�>�~+`�7�r{�vL�K`��<{�(%���j1G>�~,�#g�kuw�8RZ�DlC��g�����"���<���{������<�	iP�雰�h�K��o]��(,N�/��r���boy�hy�
�������~���+*�6⏃�!��x8�|�j���$3�W$Yug�ӟs�Sj#:�
+��3�W�}����7x����U.��Я(έ���(�י}0�~.�\�:j��D�cl�T��g���Z�:��wv���͵����T�� t�1�T4i�)ϥP��\7<l�K��7�@L-[��":�{ұ؉�<���!gώE� �`'y4��/w�EDx�.�� %Gx����L���"�B�w�ғً�I���7h@1�#��K��;&�H=ç���h��m��uQ��)~�g����l�y�`�}��3~��s� �Վ���y9��)���3羍��g���j�q�q��G�F�H��M���!�RwM>�xfNsbQB���rBfW�l�a�5����	�F#���pP)��i3 ���Zq���	�N!i���H�ګ�I�⭪�>��nވMR;_������O�ހwY����Y���۾�����6�ѱi�$
N*.{���Fd�A�hLz�L���e��o#��@ �";#1.�V0y�t~��H}H�O,
�U�Mr�TFVx<����Fp�Fh��nz�SU��<�M����
\n�F�$s/�����t���^�q�fs����q�S��y�9��i�0yQ��b�f��y����".�?C�m���E� ٥i+�e\u�%g����l���-Ҽ5�J�/cA���lrQE	�l������"��͠k���:�E�[��B���S�˙ȵ�_M�T�Z�#m,�̡/C��K 9�9�:���x~?Q�4<��-�ޮ��Y��%�s�� ��K�8�?R�<Y՟32p�Ѵ6GKAr�h���Sj�IU_cM���<��<�c�R��0( O9�n�Ӏg�>���� lX񀫈����h�h�&���To�w,���݄-�]�zd�FV���M<���i��&�2���ܢ����|bI#^zAێnZ�3R�� m����7uH�ጦT|w/�KRg߅J�D��-��� p�ƑI�v}�|v��cV<9%�^�Z�~���p U�\�h��i ����l�!�5� ����Ak{��L�Ȥ�����?%����arR��j�?C�M�.̵�ܷ,n)"]Z?��LT��](u[iX�4)�Q�{7�s�w��ٞ	��y��5n�
�� ��?��~�˯B/���&:Wi�Ȗi��d�(�_6�y���td��B�ޯ��}d� 2ۅ>Nx W(����T`A�{GU5�G��6�{�bV�f����.=��L��5�f�9&X$Μ�43^�`�pI��ꐳ���s����iO��o
Q�J�B8۵���7�UP�SDO8��3k��_��8j'���{du����M;aa�8�e��:�(�B�l
��pX c����_��~��}��j�1�v鑡��N��)V�j��
��u{�u]pC{��#洳Tf>u��ԕ�����g��S"@^�L��R�]3��k�ڡEl�/���F���9�ȥ� ��b_4_�$o�� ��v�D6�lh-�>^C�$���,���c��g�NZpK���D	M��������v�A��(�3 i*�c�h.�W�3X꾾�UHt������Pv}8#�HL����R$N��`�3�C�̽6?��v5ǹ���/���o7N/!�+��w�T+ߍ���]Rq-%�,3_.. }��V�c��Rts�ks�T�y%����|\���OW���啮����Z��F��)73�`�~��my�cO�ߴ�����	��ڊ,b/C��@n7�(2�㰳ɦ�4�n��n�2"嵰�σ���Y��+�5�J�
��*�~�J�$GEMe��� )ǹ������0����ci���s�L��vיׅp��ka�����xQq6�M�-T�n�t��E��.Ǫ�����N�Ӿ���#�O��gR���`�w�,���|	AP���Jĕ������	�����^��Ȋؘ�~Cs���Q��B�uXMC�y��}8��¥��8��#u����sM���U�|⛴48�T�w�)y�;uJ9�"�E熵�>'DI$��QĜ�Li���M�?��[3d��ˋ��^����Lݶ>$~�W��$�c�	|`uI��w�n��F��ӕ���!�������d�ݹ���'���gp��6�5��ӟ+0����Eܶݲ���/���5o��A���J�ػ��
�24��^���0��� !��k���Y�9?u��m���uCCF�{�cP7�*����ɮ�$ዷQ��U���{/������������i�ٕ��[�����٩�^ܪ������;)+o��g�O�L�Gǻ�`J����J	Ōb�x��i�5=��A�x�Zx��}Sv�:�M�:^�W1SQn)���#��X�H*6[���g�q��f��^���-�)��zF��&OĠ��n0�i�WRc���Ƀ1Ф��W�koH)ae�b��~��&a��`�|%J����r��Er�M��n�!���6���g����FRQ� M3_�o`O�.��^�YfX�7�k7���?���c�����z[��b\-a�=:(��9�Ew闎�x�ӎ�V-��w2y���{Rˬ�[?��|���~����n֞{N���!�t�P-V��g��Z'������[���0r�YGV�iXf}l:���i�@,�7�͌��F9�T6g�y��\��6�E�3��}2��<F�� v�� D���"$�C��)^ވrsHW�%�<�)竵��BP��(��n����(�[��`�Hh�"��H�2ΆfT3�J"ŉ�11�Bu�ד����9}��~;���G�o�ޠ�OU�϶ڨ���F�Ym�6.�1S躓r��VF�F�/h�d���z�Z����DLc<����vO�L�i��S�Q5�/i��m�zd�"�ܴ}����XƇ��������'8,�7
irc<�g��q���J��B��`%q!��ҕ�7 kˡ��]��'��V���H{��kˤ���0qM㖆9vގ���Z��]r#�:n�� ���oi�q��+Uu2`G��r�
�-����\
M�XR�I��#�up�{�Pl�갇�f@	t�o3�> -�a)^lB����Ǌo�T�.6�jW�[t�����t���3W9��6��<@��j���K���"`�F�}���d�?������NA�������DlQ˜�������R���e����O9Z��"b$��W_W��UqMD��,i5h�I������d��9�G;�j>.�<��~@FR��
�G�����>Կ�t�z*����� �W�)AE �%
��7�����^�#��Q����V��Z���4�
�G�l5����F�=���B����r�ߌQwtw�~����L��J��w�3����ހ��Z��Gw7���2G�o��c'��F��Ɩ���ml�B>�u!'�fīT"�:;0V��C�� ~�V�+��I��N&򝐬5�����z�c�2EտI�x����`���10�Sz	?�v���L��@�yH?1�g��2�l���p�՞JJ�(�	��~3j���Jc:��W�H�I�V�R��w��"c��o�B��i$^Ro�p���ig#��E�=��)GF���Y���SX�+TE�p�d=+eIV+�_z�0�%B���_�:L3�\�W�,j!��i)ԛJ	f�����cƪ7n�=A��	�Ԯ�����-�*�~'����]UZ�JKݖ��Po���M-�8K��^϶� �6p�؇L|c��Ī՜��&��=u��wb������U�7h윮�fl�D��1�1�WJW�3q? (y6>��:1Bi��$r��2��5��"/1=ʣN�ۘ�Gi5��=�dh�q+6�7Xn����Y�W��4|�'�4��LI-��9z^�ګ#�M-�����AiR)��~qZB-��HI�[J枘��#�ŧ8��`/�D3b˅S�wÕ����4���T���{
vH���͊���d��
s�Ȅ��7��!��\	��h��.w@�?Τږ�g��}h�0CW��J��*=c3�ɺ�d�[��]��*X���iR��k�!�]��+�s�$�:%pkJLY��ٖ�f�$��xV ?z�����:��2t�[`��p[�،:�z��c��Uܳ���.���YK�@�Z����~� I�E�T�.s)�C�&�HmQ,��7̗����4�S��ϯ	6�MVTa����d9�@ɍD	bR)Q�z�Br�Cd��?##�`O �Uz��;H�Z�q��2���G�,�7M��Q���x��Є_�`A�����0n��V�p2��Nʜ���o�u����,W�}Xk-,7�����J��(�a���L��'Ot���qE,�0�؏�����{�zp�5���,�R �5�<_�h���\"�.��CY��v��ۣ&旌������	���+�����4ݪ��zA��oAN��G���C�_�c_s u2c�K�i�m�o�c�4#ɒ�(�!k� f��{���猪[���@E����PQ�wrP-<����&�}E*-duj�'s�e�M���������0@my�(�d�Z�d�;؍/�Uj��	�������m�X�#�Q�ҬO�V������_���xdk����e�
�eKwxy����5|*N^��D�S�+�(ʦ��ZF�r;r�lH⾬�?!��d���	s�RJ` �߻<��C!�����A��q5Դ��p��aлMٟ̘�!�L��v���"���G&����9S��֝�١����Wʃ��\�x�e�����)�Q"\��]	W�k�/F�?h��#�[+����E���r�����E��E+S��^v�v^ ����h���tՏ��y��s�����b�U���[�u����1�;;���WJ�>� v�y��6Z">����q��"	�7ǱX�p�)1�bⲚs�$�쒟���lI����7�>�pYږϹ�K�D�`�+;��SvF�b�i�gk�i�sà%�"����i_�������dtw	�xtf������Z��:'wM�+���t�U%x����>$�l�S�d<d���*���_h��+����
�sS�_P��j�`OL򄑱��ܭ�Y��keg�`�Έ��j���3�'"S���¦m'�|~�%�J�b2}_Y�؝�hw���v��@ax�%,�U� �<��U쏆�kG=��q˳��7�i8Y�O	HXTbZg�d�*vR�I����lR��oo�g�E�n�T��%62�0��s�E�s3K*6�(T�t��d��tZ�en�_O1t��[�l)��t��&D�0���B'+����!)�Ëvf�C�'9�afI�̂��g��t�?�ī? ��D�
�Z��R9��?j���h�5�4�����qz/�q�����Dݩ\�bt�*b��~L"�7�Al6g�N�)� ���;B�#5�	�C-r��.�ڪ�ł��9�x�`�2������[(��|谅K.�����<>~f��O�rI��`"/����&�\I�&��6S����ij�p$�-��2��ɴ�˚��D9��o����F��k24[�P�~+�d��)�U��p��U�݈���;�%���A�0~�*�N3�(7��E�����Sqi��9�Y%)u<H"��V;>�z��5�U|u"���� �G\8������R�"
Z�NW�$�OUj7���P�
�}E{� ��R��B�
Ϧ
Y��{V;u������VpB��Grs���8!xNz!{��������(��%� F��MQX��B����0�[�kV�k���L�&G��,0�*vXt�Ҿ�s6���$�=��2��=�ڀ�z4�%��M��-ǲߟm�(s����<SD�b�Rk�������]|�D��LaSs�kԋ"��A��
�\hf�R6͙&oE�Q4r�r-ki�}�[��'~��$�� p�|��DlR{��F�Fa��xW#�<�A��p.ߚ.�7Ij��S$�!5���󦞨qcruUYn�fA?۠��n����ȏ�S!�y	e㴝����x�%�.����G̘-G���X~�G�H<d�&W?}��?]��B�ɇ�(�(�:5�Rj&�X������z��wnV���)`f�2�]��˝��3�'�̨ڗ��۩	ӧ�5�Trkֵ�.Z����G�`aFp�1��0�D3Fɳ���c�<���tHc�j��y��oN����hw�D�KF���jL/�6p�����J����I��٠HV����-W&����zZOl�Xb���L�u��K�<k�Z'�Y���f�?�-���Pn{ر��#Yz��ԁ�b�� ��*�s�azy����ź�`V���w�������?�:D�p��gv?0��3^�|!.�;�@�ZNt����6$�ԡ`=�� �1݀N,�������7�������7k;��&�s����iVn�l٧x��Au��_��!Q�t��r��f=���.��Ү�9�+V&I��Y@��Ri�D� w #>�\��@ҳ��^��W}��w��w�L/� KK=�l��9���q�al�>�RS�����;��H-��$��A�������%�NT��u������a;���\G����~��B�d������f�0¶ǥ���$�n���+Aa@2���G��`/�2-������S��<��	N׬2g�d��� ��1ȣm��a堮�0]W�V�Z���K-����H�U�y_��?��aZ�Aa\�kr���b�ܸ��Ĕ&iK-	۾�Bݟ_�T��>�ؘe�M��#1�d���_1�zφ���� ]m���x�(�~�v�7`!��������85��˲I��s(
ч{<:�N��,��]��/�EcvۼѼ8�)��'�kyBxO�t��̝�V㢝�e-�0x�s�i˄� �*���њR*Oؠn3�j���U�o��?l�j4�Z�D=40G��!�O3'�!!���u�q_�"��)-�׳��Ρ�6&K}��}��j6\��E!;�����!�5�շ1�a<His�^�^�Foe_�\og��� ݇��;�	1C��_̈́��'���1,�D��>�_��_����lK_�+���	}�
#w�nI�
��Zc����/�p��t_��y��*��"�<��)��g��!3�	��E�Y��ڱ�ǒ�r��D`n�yp��3R��dGrL��O��7ǥ���Xɮ���Ow>�.�����1:]��1 ��+oJ/���Ia���UQ�ߊ��ew�
ុ n�K� a�%HE!Z��T�0��;�(�驉?���X�)�qR�|d4�Ёb��%�j�:��9��HY����.�t�B�M Z��2<�ܬ:Y@�X@����l��ܿRm��=�ʾ����Z?1��oX�8�9��39rN��G���&诹2
M���2u;u�T.��Y�>lJ�'�(�i��(����t���ײ�u8PS-p�U���P�S����]�5�r�3�w/�ߕ{˪bc��](Av���v5���`�m��FX��B�8�d�s��Ю��߸�H��>h�'���b[�X���!l!��j�0渳d��.�1Ҡ0񪩗��;�ZD�u�g�l��DB��ER���3.X������^�01)�e]\9,��2�L�p�k(�>���Qa�*Gx�9Z�N��>��wǦ���>�i0���|.�U\���L���9�S$Z��";�z���C����Ɵ�d��jB��)���΅�Mo��^��4�&j�D�o�l������������>�I��G��l��n}�_�$�g֚q�ӭ>�"�{<��r��A��XBh��l�U�&h�� v:�����a�t�p�*�NW��ʯ֫:�]8--aD�WA�1��+�������a�����wOS� mA���}-�J�&R���2��z2g�^�x����i��(�x��C{
d�:��zQ :�Eqe����O�����{o^�T��\H&T���:���%G���˿,u���Y�e��&�z\$���W�bE��*Y-l#�ٟ����]���aZ�nC��Z"!4<_C��a����f����r�1�c�������L�x�J�+1Ā{�X @p��-ϊ$K qoa�/g~����+����X�{��^����I-8���`�;Yb�e��ݸ�`�/�x�OZݙ�e�[Ր�ڂ?w��I�V�
�L1�<��V����v�S0�Ӡ�~ѴAϪ(�j0n�_�u6WM@�%�i�������\�~"D�=b���k 6�[D9��AKx����c�YO�q+���I�W�G� y0}�F�����+�t,��m���(wP�^����Cݎ�7�@%EҨ�7#��lk�$r���
 �Ǐd}Z"�8UvHݠ'���<�]���M-�$#C�C��ƈ/{�iY �P�.7����C�+�f�zm
,��.nnPC-���g�Y����dm��7}�x�5w�U�Jcq�#�2��>�b	J��b���XFq�a��8��V�)%X��8bc{|�C�ϋ��ʯ�D��f<�p��hv�xU���/�m]]_��V�/��A(=޿C3;��B�%k��(S������Ĕ��7��Sޜח/��5yB:���z/�T�a��I�w��)	O�=I0�s��&� �� W����r���`�
�����!�k^�_!����qJ;G(��W�$��;��Z��,o�m"ƅ݃�*��F��G�J<��/�F���Mu�?X�v�����OB_��f�H���^���Ov�ǖ�e"�V�k-�4b뿄����{�'#�������88g|���\�H}��1n^	�:}ؽO l]��
#��Hu}Ǹ~����{�F"�4ީ�m`����I�=G�|�dA{�#��#���$��C��%�Ů=�)>��A���jE�%��~��zw�q�,�hפ�Ơ_����UE���Ӛ:��n�T���c���OGySK���}��n��PSl�����fJp񹕬�X	�;K���f!��3l�@�?9�I��X�E�y��S��D���{��_~L;���ف�v)������J뒿���f$I��r[s,K�t%����̞꬜=j�P_��`{C�+���dy�!�0�׼�6'��\�\y�Ko[:*�vv�I#9e����R�G:��RuXڸ;��kU��� !{����ξ�sʛ���j����G`gM(�H{5b������8��M	�Ō�O��r����e�k�Nes�V�w#�6�������넏�;��������m'���ZF�`��\VH��l�M7Ͷl����42��n����ޮ|��)��f�n�d�w\g��k����L���03�.�A��cdb� �cM�)X��m��&%��ȏųy��l�h����|��4���z�+ +���R-�W@��a��EP�]�m�;oL�˰�'��u�	g�C�9K�'�zu+c�>�����z��Ø<�Jm�/�����s8g&d0�z���ޖ�r,u�?�����X�rKP����8��ł�Rs)��ū�7��Gx�:�&�Xc�Ԇ6L�����I���.�嶢d�8�mۉ�O���y��U�ku+��\Tg+4U.��n�&v�<W�9k��4�I�B��t�������my+�@�N�H��5^�\4�
p�}[?T��1��l���w�5���\A=��e�mM޾�>^�)�7܌����KP�vYɺژh�����6#�ٲ�o ���_ÅE�ЂS_��%R�2m��z]-7zS6S\����T� w8���Cr�t������V�O�'�)� r�Qn��x�wMGs�8}��7#eD��R�%�a�R��	�g�#'�)�!{�,Ox�g��E���?S�Bc56��<o�Z��!�Ռ�p9O	f������Uj>A�q#gxf��v�@x��~�B.�t=�W��
L���Y6����'�gEqehxW9��!:{�Rr,��x���P�b��������+2�nH���i��Ɖ���Z�6�|?:�6�����e?~e��l�d3:�Ts�
� �V�Dz�˹�m| �&2�^���4�΀å��ٮ�|/֭�܏���b�:uD)�Fj;���A�SE�${:jCe�%�ҋl�p�P 4�A��{��a}^�����R0l�f�t
�����m��d6�7�:r#�iS�M�{�=2&ǆ5�v(Fy�W�֣	Tӿ���[F5�(Y�/����s)��D�f/2�9�c|8�Sm���XK����h����ߘM(t>�|լ@���pU��.��u�rcS��o8&�N9���'3�������o1�v���儈'7Y�`�^GYa[�6e'?oO>h�No�J2Z/�+�o�K�LS� ��f�=;j�?�`�^�f��H�8�d��&��hdh��!�eZn��#2ӕK�|/��Q�����DK
��]�:�@�9ƿ݌��sd� �|�<wd�,�p����F5�Ib��a&�݀N���7��^�ՙ��n`}��脟^�yo��� "���u<�J�#�.K/@w��D��E���9�ޔ���#�6�
��	$N%�ipZ���[hP��E_��
b��R�ˀW��کUG�^�C&�l[�.́'%:r�s �XAW��l;JI�� T�9Gp͓7T[ː�⧕�,�
M\V���q��kEW�3n��(QKq�M����y9�R�u�W��dH�6Dо��#�ݖOIQ
�ў�y�TtmW�H9.�E
�w	�.� x>��	�Y��l۰����[�p,? �������r�A�I��!q�39�/�7�cᜆ����Z���"u��.,����ZP�)�c�
ܻ������d�9��>~;�U�$��<:k�e�_/it���?	���'�EG�gd�t� ����O�k�^���t=}����Jޓh�XkG�R��?��]� ������	%M�K�2��}�7��MZ��+�#gVĶ��~1�Z�J]�J�!�Z�	�y�K˒����>����cD�>m���NA2�tޏ�s��2
$JP����4Z�p��U#��=�v��Rh�-�
��!Ln\���|���K"�m���f���u�>7��9@��=ΐ`��t�H,�f����%�p�E9~���s�x"`��I��KB�(:IL���;�+����p��!̀�]� �,�V[x�~/��O�����'bD��8A���$I�/�U�o}݄����a�38���5ܗ�e����P�Pj�Z)I����_��,@�0��t7�
}�_J!hmJ��A
�p�J��'#�1�<z`�!	�Q\*��� ׽�����p���Eo�Qp��B���4<��Sp���zy��+�s���) �;+B*$G��O:\=�dnT]�UiSj���6�U~¿�2:b�d��TR�)������q��k���dTH?�!w�Di�B�Ð|�o�_�y�:���q�Q.�U�@�(m,@~�ʠ�<t� �OG�I(�['���W��uA��oY���Ͽfr�䩓�`�E4��e~�$=��*�s�|�Z�<����*l�E���W&Nre�>�&�=
��:�{��M!%ن�̮�,�
(W�F�}Y�)T�b������@��Έt!\�]D�����iv��i�������^�����}q*d)���O����[ �'�:)����y�̥D�Eq s��X�x��6Uš�C�;��a�s�e'�Jl�[y
c��,��)�m�� �'��'4���u#�2��p��~	n���K1xP�W��t�[��V)��"�9n��F��i+��svK��i��*��������%2���%���<�*y�ȡ'�1n�HD�U6������+!�!��-=�z�.cP�Ta�Yv":���Ww!�]���?�$_�g�r�5j��@1��wEh���wʡ�[�+=��1/�ڼ#����Khc�(2�l'�䮲�)�&��D�C=�p����զ&Q�d�ғJ���c�%daŊ�#C0{���{BUZ��ӊ"jSj�����D�L].�ټ���1_��z��!t��+w����b�pl�CK��uZ��}���P�塙��ʥا0|z����0�h�����d�H���ܪ�|�IQyd<�v�F��^l��9�/l�/�HH�1�?4m�YӢc٣�ߨ���Y}���vh�M��JJ�0?�,6�+����6Y��ww*>c����^v��r(2���W�d
���b�,�i@�!Bks�W�y3�s�s��yaC����^���V�����}�e�+���l<	
���A ����@hS�E�o˛��싉ƞ�Q��E��s�[UX�7���e�>Ӏ��~�w���.N�L �~��0�h�*�e�BJ0�e#[��i�g,�n0j3,|��Jct��vr����mt�/dXg�q`ή)�0�$ƲP�)�`@��]AL6�=�w��:/6�1V_�{����` a;4�v(V.�>�!�b ��� y����z6��[�,:ߤ1��U�$��y�I���DHi]Z
�o�q��wM�g؞fzSY~=��\
P�,>L� ��=S�.�w1��}��M��
3��x�U����$�.�;KR�̫>N:�z���P�
�WW�e"���@��~���!!�]���F��K����3[*łF�Gۺ"�2[͂T@�����x���LJ���-+N{T:���,ǵ�(v���Y"A��Ee��CP���]'�~��uU��A��3lr��'�ǻ��"�M����A�i�/&���2�����*7�<���k�k���/Q��q��B��!��d�}��^�fH�L�_F�}`6���Hh�e����XW�֓�.sd?vi������	?rMT�8E�w��W$�`+r���}��c�l��qb8�74���b�2GQ�#yTJP ZT�VL���Rb�%V :�s�����R�?��<
�_����T�?�.]�[���lqC;d����xk�r+�]�7ͳ�YA*��ζ֗���\�1uh\c'\�bq����ܓf(�،_�Y%��9��V�e��|����l��#15��M�ɖ,c�??��-C�.��
�-y�UN�7���h��&�R$-�s��ĹT̾r����
Mma��V���%'i�(�J���؂�����߷�K���G/���w��:���'�F�#	�K���rH{ڻ,���k���������RH�����ߒ��n��*��k������[n��b�+���8p�ԭR�����=��xa�xY�Y�$b{I�Q1���%R�2&���&V:�Dd�]P�P��T]婈I��XC�V�a�v�Ǳ6�Ě#����"�X���	�	apX�n����sf�s�:��i�q��%Ę���z����\:��zJO{�C�r|fڞ��!�E�o����I�(cty�4�W�����r'�����+�z��� �[�e
�0ZˇM��+�����o�9;��rz����3�%����kц��bw;��G~�����@8�Rw�ˉ�̝-u�@-v�s2NU��XWS�����&C���ο�yه��=ڤ�(�W =���$o�[�3�Zp�1�*�س���12�����|_��(�<sMة���U堵E[5���e���z�y{ �O6H����S�2�M��0�_oan�[�֨C�����#�u=�Oe5����=�&���#EvyM��xt����Ǡ-\�~\��76^�
��Z�������|�C�2!�W}u�� `�P7s$�����]E�ǧ;�7�<όKǄN�m(��'{-�h�qRo�#|0��ղ�^�tB�Ͳ�[���Wό%�b>��d-c(БU ��67_P�(*��<}�����q?��k�Y.�ᰖw��|���0�s�Q�l��?��4�ԝ��Q���[�����}���7;�k��k��0�Xӓc��� ��
���"6�y��֮:1��e9°9�{.���S�Kz�$�Z�P���o�_�jbu��ϿaA����w�>{�����
�nW�^��f�k�w��+
tdl���&>�� mۀAWZ�ιf�{��p](�~��vZ�����Y[��Hc/u�&"��G�M���nw�E��h�6
�ͣ�+�@�t��v�e[m� �Y��ݽ�9�L�6L�}H�[L����`��2�!S�c���A9�������ci��+*f��X�5�0}<H���X ���
W��_���ǰ�D2�`|���Md� ��$B�k��ұi#Ȓ;�Du��̙:����^��;���A��g����-������<� /{����2f�?�\X���^��G;��fᲧ|m�j��ɢ�K��I�Iǝ�x�$�2�g�rM;��\�v͌p;��z������R��Ju�-s^Gd9k�
R�"B����zw��F��\[<a��1fH�����-Ѭk��C6`��e<a�3>��3���hZZλ���{ϹOê����D��4��K��dl@מ��"o>����[�� w���vBA&��[��m$��uv�K"Geލ��&1���D���1J�I=6�(ͱ��9�$�N�N�R}l��13ӂ����ɾ�8��0D:U�)Ƙ��:2�q�=p�-�e�A�7���K!H�.��?P��v�$Qℨ�5Ud�h��OSrNV�tV5L�fg�N�蔪�4�w?���ጏ�&�����QQ��;i&���>�'�B���bY�i1|�z���]�an����b��q)�[�T��
������:���yV��Q��	9��7�:��6VA����>а��
�]U5^L~ɦ����XI�B.�j��,�����Y�#��G�i��ʒ�&_��T>����S�ǳN�4������S?Pa$��P
|,W�u���ׇ�w+�m�4s&uM��զ�z�r����h`E�o��Cn�h����A�������Hse��m_�g�zi;��� �э����K�-�U?�F�A��=��7�$����Zet� ��/��n�{A�-<\[ߺ���.e�9 t��h8Wӌ�������I�m�D;��ob.�s{H+�W]�$U�Z�3}_n�1�/u��m�����m��\Z�-��mco�\r�>߄�|����ZNYxx�Q�f)Ϳ���%�2���[�t�$���?����u���*x��
�<vS8rT�)�:�����=]f�5���|
�áe���䬼}����w~��}��Qs�M��d�c=$��m�Oo��
�Qo����L?�c8�`��q1�{����%K������$��Aj��$Ԑh�L�$�֢K�]�+�+5d�tXl�IV~�QWdr@��(����kGZ��.����{gq6-����쯢A}Ê}s�s �Eܠ5VJ����uv�ߡB�ΟإCX�-���_�fN�=^QE�0��|>9�}�÷̧����e�l��%e�W	{�)`D��g�|��orIƟ��Պx�/��e���3;Sn8�K
��q��YB��p Ĵ&6��J�+�AD'ؙʡ�oE��|X�qj�vW��7���n%�1{���D>��a��8<���֐�7��v���Ia���k��K|����r��SŬ���t�x�c�%���[��eo�h��*���A`T��� d7����ƶ�ɡW�v^�#��`��"�tD8��-G K�Q7����#��7�j8���7ez�X,�z �}
��Ğmy��>�sy��"�M4^'7i;Q�R�.��@Lhc�~lz�y�u�?���MZw�w�e�	}ɩ0�z�z��</�׉RG���'J���1�_�6�Y�[8P,��ܷ�*�^v�"���:ک z$p�>�o�C�)�%}vkˈ	���V��F_����@/��l2��3��k�}��L�XH��� ���+�>�V�ӹ��F�UY/'�|"��X����D����%hj�`��f���,��G�8O;�&���-�q�Pkf1�.�^ghk�)�|@!�G�	��Dw���C���N�MwS����j�\&A�{���<F� �R�r�{�Kr�`��.���ղ�h��������-�!���NϠ��B�e)��ߋI���Q�("���NF�[��1FA�54�νH0�' �����失��9]`����y�q�TJ��N���]���G)��*�����Κ��2��L��qNPR��C�]�'��om��u|ƚ�y�+�j���5+e*,�3�b^�r3��C9������D����^h��$�޺�ݬ�����t�󧭆:/��X� '�;zp�ɓ��[���\�ڎþ�Ϥ۟�G��1n�	]�V6� `�G���w���6>E���u��AzF�M�Uw�=���U����f�-xD��u/�L��	�	(�en(2��{:�O}�R�f0�C�����8��9�X��X��`³�����fK�&]MI�T@���`U�fo�)Ń%����S�a|〞F:ZS�����}RͦQ-	h�T��m�)�] ���B��2��p>+�;���E_��@<,N�}��^�I=��]yÇ�E�L8�)��Q\/���C=��FD�������YG�k��/_ֽp�C�!1 Iʪ�������5�Qy��2�P�F����$�D���*3.5U힧��-��`yb� �1�e�2R���؋�~A?,&.�O';hlP<F�7T$О�BE"a7�Mbp���Tmp��@y�'��x�^�̧�����"��������,p+�=�oW�冁��@"=O�>|��˒�������q�\��&gn|���y�՚2�b�ڋ�j>�Ǧ|����ٜ����*�����oD�	ؼ����:�c�Kڜ.va�0�gz�}j<��%�
!O�]\h�dwj{��,���&X8h[_Iԙʰo���_�V��5�Ȫ������yb$�Dq�I��i���!��u����[W�d�;�U��'!bp�āD�\��_��	�k8^.����A4��:����']��3����TN0%�ܵ�b1�F���8τ�JE^b�I��~a�(N���n��@^y�sՂ~�p�����Q9�5���j�Yy��[񤛈��0G��D��Y��x����q�$&"���K6'��  9�;��%��S<�J�}����u.Ni�p{���;�IL����m��������r�ǻ��F�u�?M��~Ԅ^��s8=g:�e�,��$��X�g�;�'R^�х�eE���,K����LA�v�v�Ob���z#j��-+��Ĩ�!�߱��2�_էk%�#/�ť��_�|NJ��0�<虸��'$%��):-!�9&�s=P)q9�.O)Oڣ_�U�:y��ˑ}�
����gI��'3�=��)�ɼ��q�u, g"�`	�;��'bPRTO�j�W4zy �>����UARD��0أ�!�~�x�0�(!�M�qoR3Ds�a�W��ۉ��)��Z
T�0 ����k.����@�H�[�z�l)-V
RE3@�!G�x(vöK���$)�vM����t���ٓnXʬ��2�!�H�Gs2e`�[N.��R��X��g��G�ެs�o��|yܓ�Q�I��(�"GFɺ�E+����NɼFWL��Q�G���a�k��%�]���RHYtX�̗���k9{�=��O�8�-/��z�SI��O��Y�@H�=V	1EC&A�K��K�1fI��oZ~	�S]���y�A��&��e�UwS\��+�4W �E���[m���œc���אGt4T1���v�lML�U��������iT/��x��KM�\R�������N��F�;j�Y�����>�^dy 
i����L"u�i`6}��L-��m�H��/X��������>���Brf|��L�+`lLc�}�ُ3����d�hV R����@�`Nq'��)R����{�����]���1��՜�f�z�4�e-�e��aL	�h!B1.�֒Mj��(�A���9\���fB=K>����y{�e�8>w��֙��^4��u��}�6[WaU��ie�a�]��Q_w��_`�g�`a�������R9�<�G<�_�a�)�k�ZF�������b�A��}�K<�6�4�E&v��>�/q��i5���M+�Y�׮P�#��:���̸����D�z1b(b|G���l���h'����,N�ȅ9�W�W�^A9-�Li�Z��6=/"-�Yп:P��_��f,��ȉ�rO8/�hA }��k
�
�jgL�����^��\ԡ?�����_�7�JW��k�&���it+ar:T�L�k�����7�_�L�~j`+p��~C��?�#u���q6�����!	�/�M\%LO�ظ.1��)yD���a�H�p���ӛ��-�'����]Cw��u�sv�,�%�Ԟ��fJ�b�#>��w%�=��z�\F@I#yD)�3驢������T0�+.���+*w@�"3������;�Mf�:�D&��T�k�A�a��b���R��)f�Z��dj�&T3}7�/��>�`6�+S���n����|��j��&͚���r����6�|w/͐+���H��7N@壥��cS���@T���{���g��_X���=?�aM�fTZ7(!�W\欭s�%�|>����92N�۸�dH��*�,��i�(�m������tI"�Cn�����������G����\_���42�����*T_!��]�������d&B�1QUP0�m��R�͛٠�tU�O�+�\%=X2�1>`��#$߻#��8G׀���٨���;�KZ���zs ~��+z�>&�{}^a��猺�o�	ңܕ���?��y��4���@`�k�(�z�u�(�A�W�s�74k��D���b�G�@��EG��]�s� D�p���D��pn�E���d���M���=���숀]���G��a��Y4��e-L�. yY���������x�՟
�gdh���d�<�H�E��%�����vE�z�3ɄΥg��M? �o�(j|B@���y�}�濋 ���=4�-��o k?;.C�ʚQ�/�` |ja��"%O�XΖ9q-�2e�_ρ�`���n�}�cn/�G~Ր�j��M�w��̇qyP�B�����ap�s��������m@�;�<^���N��'�zW�׶����޻����z�:����D���i���`#{�f�ʨ�t�ާ�S�rz���_�dYAo�F���n�B��:����~;I߇��1/��3�L�[���q�Bs���w��K�E��[VbҼ�u�����\ �8=<����֐�?r{��{����H�7�&�<ݮU����Q�Ouh�#����8^��Ƶ�h�� ��
\�Sމ!`�x�g"�(�W����:�O��%b�\Ǿ�*N�c��5"aqJ� y,BĮ˘��B�M�|���>�����f�3D������B0��洽%p؄.����cIbG��N?��N�o��I*��(f��c"x4T�j�
"l^�ͧ�<���3��*��Az�E�i���V����E�3X�����nWs���XY6c,:���K����H��E2���7�!��n�A0�QK�3W�������e��u+o�.v,{g��K[�g��4�̛�^�3�V��Y�{�0$y]�>�Hmd��p��iX�K&a�6{�<N{�!_��ū�{v~�G���FxG�i�qfy��� �1=�l.Ȃ+/*�[�	���`����G�=�4��
@�~��|���}xJ�6W-�(We���G������1x#+��c&��ڝ|@&�!�!�r��?J׹�V�G�u��:RP6�d�s�@�9���v����w� ���y���|�y�Ͽ2�T���gn��z<������J��?r+uk��V��r�����ҖGk�w�+�c��8
�b�
a�ƒ
�u,��/os�I�;f0����I��Y��1^�tD6�B�W�?׀����f�H^&H��ޏQ��zB�wȣ��1B���xU`�\�qF�O7U��Ŀ��(@�L ?���6��Q�o&�ԏ�ݴo��y_!��ő����E}O��Q�w����D��$[3}�;ȓQS�9����wj�c���?��x)��x�lj４%L��l��N��6��+qѯe���3�6��#�-1T3�k�*���;����p�����ϸs�>��֤�r�3竅?^΃���X2��f�=�|, ѿ��9={~>0�!'ݡ1F�c!�c�z��(�%4e)����t'Q���(A�XFD�eLϴ��ܖ6Mz��3�b���D��{���r�"?@E�ި�bs��/�XRfǦg� �X�r�PW(����k�j}<�w+�؟J����FO,��B,�Y��+���W�Uq){������r�`�&��g��3F ���l��O�)ΐ9��ɧ��O�w�Xt�HA-�{�P2�~��$(b%�^�pl�����)��&����m�ϵ�20�~?�[h
߷���9 E���-����d�e,3ޕ�_��U�ϛ|L_�ҒSPs�����ƀ��L�޼V�� ?_j6k�G�<���j��/�I,��}ı�}��v���]uh�������䐍WS�εL�sb:7����GgƬ
��-�H��{2�B�ϒ믓��.&�9�
�a�)�㯽0+����V�$�0BR�iпB<S�����CVPP��j���`���,r1{O;�A�VN�Q�T�8X��p������L�,��(�S�U�=c���I�������U�%Qn�Ħ jC$��#�ZH��w�3�JAN��8C�x�+��#5�;;��S���Y�|�FPY;cۻ�$DP�}��x���;qH�+P)�b����2zx ���@��5�g�qC�`t�o~'�[Ƹ��?�˿>L3�a��~�'`E꽔���w��W��g�k��Tw�Q�Ԁ7�ZH�����Г�ض��q!Z����M����;@����mW@+Ȏ���+x�8 �Pnf���BEvC@Ý����lK�o5uGh�s=W����.��:�QE´\�{≎���5�Չ�0/͗�n���M�%�����˩W���	kl�T)7����*Fb7ǼPw@�3�r����	ua��R|B9y0ˉK{P��Ȟ��Mܖ���0��@5|gl�BR�mWڕbS��=]�7c�Mئ�i�"�ߨZf�Cʯ)i�<+s0�b�k�Q�A����f���J�������T���6�
�M�K|��,��d��(`f��jBH�"���`�$W.��
U��D��8�����dYkk��ɲ�C�S����cMf�{�\!|2Q��$ؑ�S�MEp�y�LQh.��3�P��w��p%y6�s^���wE�g;;gZ����xUs-d�Ѷ *P���xF�2���.q+Q��l[��0��ws�m�ީ�#F�y�l�;����r+:������'-"��]p�V�!AtոC13�5�f�H�-���D�
�f�b�w|��"*Õ�vX�������AB��dr,�^��p��c���u�m��a��gr�u�bA/�y����tI(x���zs����K>it4�`�:)��L;?GC*chr'����/l_nM
g5�vRCF9IS����zK	����������@��dr<aÙf��`8�16pwu�_�=w�y��qt�_̟���r���n�I"(����D�K쇐Iߍ��2R��0����|���G�A/�H]��h���}ȽK����6�ou�!��	�ʫ!i£0��c��liP"�����7ԢF������� r���9��e��E�e����w�0�*_et8�;�4#�����E��s���.w0�K��Ed'�K"�.*M˔3G?ue�K�Zp����%T��ɀ/��O�RGpԷ扂h��WVPM�3�H�t��p��4K�����ڂ��fǢ��e5��V�IԂъO]��\]�*�,�rU��,.agl�|��F&e�}�p��:��C��e��(xw�F�RMk	����/*����r���z�Į�n$Wu<�;֘]�?��F�dب�af���e�_{ZԐ�M�y��pl���IF��0D�V���@� l���UެNU(2�P��3�]!F�6��٬ p7g��0��O�9Y^?�������]tm�"N�k_�`�\D"6�\���]�-:?wZW��Ơ�4��\��>,C���QLwwĉ�MB"��R�E�}��D���Y���>�:�*l�î*�wQm+A@���������En��WxN���y��z��읅��	�`����(���b��_��l\���;^>qc���:�+�dM���qL�V�����TUE�ѵA>��7��/�P��r^n:W�܍%���~���"��p��;�	�(�U��[���V2����t��JV� �t�@�62��%>�`ѫ�n��)y=攞D1ӯC>��т9�ȫQo���&�L�$ب�o˽��W��� ���@	��Ր�Ҿ�H��X�������d�����"G�	rm���7��&Y.5 ��M�V~�C�(�
q��֣wٹ��BXq��yx��EuL1�Ω�f��X'G1t���2��rZ�kDpT��WI'y?g��4�/,w��W��ݥ�8k��A��e[��.1ob��M£[\Y���7tK���0\�=�.F�'I����� �ߩs:�l�$.�}(�BD���ㄴK����?;Ş^Xq�2��'�[�;E��x��%�G��)�ЕK�$�mK#��M C=ʖ˩�"�g�]�MW�v�"��k�r)��0��`w���|��	XC�;����8�t��8�����9���ޅu�d����"��^��D{������������O�m'���R�#v��Z��	��.�������Y�XHC�uҍnO׍�����B�����yS˕o�F�U(��$an�ŵ���*䥥�H݊�/��${�w-����k�5;<,�&廌S>��F�/��%�>���o�!��TrS�9�n��-���r˸����y*���"�\�0Il�/C��_Ӳ�`D�`���l�U�5��uk �%�('�����Kn�0;1��!�zr���U���k�h�a��2?�=.T�y?֪��Lp����%��B�H�?vf�q��}F�rx���
�1�-\����m�zZ�F��!��ZI����g��������s!�I7��:���:�}!�������Y�8�ƨw�6�;�( �E���ƫ�cq���*#m/?���HA��bxe�@4t��	��'��<G]q'����/�ӟ_L�,^*��m.jRvT�{��C:H��G$y!ҊW!8�Zn�}�%_�MX>#yI�V����+bN�M�`؁{�f}ߐt�cA���H�»���0b�����W(��ͯ{��q�S�A��6�iSnt�.�9@�Үڱhio	�v��}��v�2�\��W�\M��Og(t�{.�g��Wn��ԕ��>�R�gS�+�;�b��jL]_0���z@B5��h֙�ߖa��-!�`8IپEDo�����EH�)�,��T�`OӤ%��**|ݱE���C�dC�R<��=�e�yEr���N�ӺCp��EB�6O�B�&p�o��"��siV���s�"��'WW��8�~�����ߺ����KPr7���*���!ꪩ:'H�:�!&A�]���]|��J??/Kb@D�i� �X�[�B� {��#�]�m�x(2�prp
g^Pa�J��S#���ths��Re�:�l�0��zOws�~r��N���X����&P�U�-�nP˫� ֙� ���l&Y�=� ����<	|���	��k��ÜW�ڞ��߰��b4GN� h�+^-نx.G��=g
M�v :���<Oeh�O�hɤ`<�+k�I�ڨ\�D�� ��tR)�(�5�� P�Jb_�����'d���-��t�l�VU�bOT�Z�7U1\�j�:�d�U�(���}��ϗ(��+����>��� y|��4 '�C��7�OY؏����;�]���%�I�G3B�O�=#�١�8�	Ü���j>ٛ�E�s��ӫͮD�eA7�*n\�ɑ�\8��8T�f��sPH� n��kx�]����	��(oe/�My���6�x T�x	�̳r��Y�)Q��!��4�z%��j���n�#j�	�\?�\�:���h{^�?)�2a��|J���ۃF�P��4����4q�C3msx�9�xI��������ص��@V��ue��cv�+���~l�yϼ��ܼmMA4��"�U�q��b<��zØ��3�９ѱ���-�����MA	O�7���\��KY�a�v$F��6������kO�wjM�@��T����v�R\����{ ω6��k�G	��[��Jm/�R��z�R���,��1h~�<�9��䢁H���!��"q}����qHiW�ł=� s�h�\���z{��ϥ�F;�d�ꁄ��!D���^J�ov�t�����$���]��TT����)���&�c���8��������ȃ!ta�/���p��ͳ��򽓐�~�R/�Q�+�ӵ�hC�Ԟ�&g�:�J�/�*�U����+�k�nG$n��Tu��X�j�̶���ڮ1��7��3A�@uU��<�����
4z�;��K�X�1$|f"���r��~c�mp�o��(c}u ��^������a�#�;��
�v ��̯2 ���~��hIL��!sGk#-���`gc#7����GD�=�miR*S_��9��r����FE�,�9�����Y�o��2/S��@bp��԰�ŏ�a����a}�^�a� R0�zT�|��6�y��,����B��t����'%����m���aq�lHI\A�tF���޷f
�*�3H�,������mh���E�1g����Ѓ�5ys'�ޤ�P�	�E���)�\k���d�~�>)z�di�5�ɒ�6$�V%�+��z4�������n�����0��X����Oax���<���7���3���V���H���@n�e�,r��U��t�,��R�NA��|����p���\t?B����H6S�+9i`��W�)d�J�t(��P^|�	�u�2��	��8���ſ0�3b�6����2OU?
^��p���xk�w	ApE!��h�7�d]o���P��yV۬�|Ab�5��:�x0�9VS,r{B"�ԂU�"�X�iY��*��x���.a�{ @�?�
��jU��_i�A��#���:h}]����$zbM��=�!p3�U��K��#��/n>���;>��q�;R!�RǓ��V�z�<Tؙd�̬p*A��r���Q�����.�X��˭�+m���h#���;Vk��'�YMZN�pH�H������W��.\�4�_��S_��{r�8�����B
dW.��k�_1dΆ��@ݖ�^ƞ��_���Hv����q=_���'����}�Gp���;���qZrT�vZ"|�t�y'�c��	�RQ�Yaz��х���}��s*�g���`(�� -��j�܆*���h^�V�O��Yd'����P8�Z����٢ �+�������يB�'bܧ��b��������;^�s��l����Β[O��:�ď~�C�oFduGIu�T+:�f��2�<5f<̭�~��Mb��H�s:�s3k��0 z�A�z�wf���ïPcp��r�Xh�j����?ݚ.�h�\�zn��\� jԙOi��~1O�[��|�fh/��2��5/�e\(C*q�T�"���o��W�>s���=�ٵ@&�N`Æ50mR�#c���S�qȍ+��#�YFO�_���l�ƌ ��\��/�`�M�1L��)���,3l(����9��{n�o��%�}��+��C�d�OE�3���p���S��L-�O���%�
�W:�������P�DUmq�T�"~���-}��(צ�켡�[���u�jVǎ.�m{�wɘN�V@��^�
	-1
U�U�&���Ds�~JMT"YMM�ӊ$�ύ����OQ@�q`�SlK�i�����ۭz�QẮY�rH	"���/D��p��j�m�^�\�ھ\�Wκ1�s�o_g�c�_[�t�R(���Mm�<���|@���V�C�.^!�g�O�& �h�vǃ��Yy��+
��>�����#�zp���^��	��A����O�`��o@����E䯃�ֵS[F�.����bJ�j�M�&���ѧ Est���=/n��6�*dX"�����^೉à�z��	B��Py$�K$�ҷ-��pK��h���F>S����j%+#"��?BH'��E@�?�vf�@��h�w�������{mKN)pX��ҧ�������Y�v�kl�oJ nK.N�G�~�jI�4�7��������s2�]�+��h��D��Xm�u�w��`�(��RHt�;��>�f����\����f�=�+B���׍T���f�|��-}%ޠ�A1���ÖF�+Qo3~��xUY�z����;�蔺}
����q	��Ꮪ%�!cn�s��+n�������L���q~��J�{>e�;� U����Ŧ���'���j�c�P��W6ʃ��N4�+�.� O�Y���`��!�*Ʋ��vD�BJ��3��)��t�.�w%��Zp?���v���{N؉D �8K�+��ܤ�QZV��o���a�ohݮq5S�{��pzd��\�~DE>v<�׫�/̿���G (�,dJ�J/_T���{���<6�)�P�D�#ٜ}��'�aL�t�����y;�֐n0�.��$�v�6�}PUax����.M��/B�t�U�DυWCf񯩲A��R0Z��f�m�\ew�v����=K�0�k�3�{��Q#q��� �A������V���.�0��/�㋇���q(����$I�;�ȫ�nNVZ��<�& PX������u�!��('e��u�ǽ�J _`�W�Ť�=���25�ތߟX��u��M��4��{/�b�9�p�=^�4r�\3R�����(�mW�� R�.����rB�t�5EG𱒆�	h���w���V�0J�n��4���n���/9�Ʈ������rW�x;~��pW�
nw���\��~Sc�ZL�d;A������9?�21�	�*,z��`D�o�	>e!�l�aL�4��֊����)[E#���U[P<+��,{	�g�0��ߖ�:�1�j��"������x�����4L�z�c<�]J��'t��C���35��%,���
	j���{����u{y���A�쯄���G�FH#Y�ۻʧq�������+)��3��~P���~�*�D�`�鯀h�	���Zߗ���$=��%:VuTg<tv�M����u��|-��T-3L��#wt�*�x���J�0�^���bn���э
t�{�i��W�����Y����6
��h
v���E-�mi�&��`�a�!.�\�nu�i	�0���/N�����Q������e���ѤsH�ľBIMC-;VJ��o�K��j�f��\�@}e��aq�ּ��Xe��A9�W}���;߮�����r��$]k�����j��c<��ꬨ��ɔ�E����������X�z� ����B׭���f�Q4��跢A7���a�~η��?�_'��ŗ�ꢢDR��̮��vAc��F��B�P��VvnH�c��\I�t_++Ŝ�����aW���8��R:�n}5��B=��mU%P�)U�n��"9j]ƅ���11'��{4��ԦC��dq�]�S��\����p虆=)[?�Q��y#%f�� ��i�s�|(y˄DE��HӐ�̱%���}�l��^��f�eIS9�Y6�����5f�j@7ӻ#���� �^�\����c	��^+�b�3��C ����/�N8�Z����M��w�t�A�b�J
e�R�������u�%BM�w
T��b�p�Wo����R���b3Vct`� �Y���G�.���c�i�,���W�񑰶�7VX�;(-%8��w�'��<�@�T7UL"��c�/���C��ؼ�۔"�'|��o;ܥu~4.T.戊�/
��uV�	^D�2����T�=i�R^���$j�M��:���7Mp�����@>w��L��g]o��z2ꆨ�ߣ�Ͳ�X�H|v�����g��hE&����J*�����`��RU��s��qe��x���$����{��b&Q��������� xb���y��dg�e��<A@9s���ό�h�Y�1�h#�a�_�nk��U�q��������:�PNT��4�ި6��9��{��Gn���%X�j��\��P5����p��~۟�Qw����7G��{1�k��G {�h�Vy��9>v	f��������Y �0Mu��N���f_��v
>�i��̟JO�C՚�v����hؘ���e�������jVs*��^�_��xk��w;o�孎�|�x�
a[s\�=xY���z?o
H��ʲ[P[y�Q���2��tޒ@���t4�V1�ʼ�yS��� �e�C�,�JS�OF�7��f� )W���}�F[؃�r3m�\^ט�v���e(������CN�_���@j~�x��!�jUe�9fce������w��)�L���FP�����G9~��p�pV794�A��7������E��i�v����*�����o�b�#8+̤l�B`��hq�C�	(�S�?�ȸs9�n�e�ާ���w�u�8��ad9�tP�����k\
U����pq�7B�����E*����ou2 gCu���7`�op'�Е`��iʨ�P!���NvPY&������ i<q�h��1��n�5p�X+I,Y�)�'�A�;{�i�@��}�E�6ʝ� g����� ���H���?M{��;�P��C[����9ǡE�Fr�Ι.��>�f�b��l��7iX�1;'H�:i
#g��h��u�6�+�既p?t���S�����~��K��� �ƶ�8�'�\���_꺎ZX��I��(�}o�sw�t��d�G��k� E����DJ��>��O�7��|���
���2��wSg��`[Q�*9 ��{^��Oc�{#+�s��S*�:�Q@z?W�y)��{�q�7Sy0�-B�y�>G.��ӱ�H��;x�9�o�f����� T%�W�`�3ұ@�x��G�\��9�$�_���DU�x�6`y�(�8�t�F����J���^���A��7��6�t���/���y��Ƹ9���n�R�:�:�_�͋
q�{Y�)����p�G4�m��R>L��`��%�>p��9�Q��C:V�l��[�,k��>�T:6o�K���ۮ6$^쨬ŭ��B�扵
�y�-�A�3FtD���.�"����\ !��d�F�/���um1$E�{F�Wm�>���2�[d�q?蝨����`ؾɨ[��=`���XU��U��maHR0�]� 0��\)����j<N��X=!�8A4-��{�I���<t:�L~E7R���3���&X����7܅�]�V�D�	�޸�q��!�ݏ-�<ˤ}yC�uQ(����bt��N[=�H�5���`�?�*o��&�d�h�PoA�*l�Z��ò��r�ۛv��K��/����In���v�A/Kc(|3�k�`1����==P�O
��Ôv�@e�"[|q��H�(�ܷ±:�,���(8�6��-ʪ��F�c���!��%3*ڄAԤ�3[���K}�`��4�V�<1��Z"����$^���B�<\lU��ng"g�j�ȉK?_�t���X�_Qd�}!MP|�x�D��e����M�/�@�i�!z���tt}�� ���	p=�1x(�D�[��U����� ��I�� �c���ڜ�A�.(����YӪ�<[�>	�N��3�sV٠h���~�
&
s^)b�+�ʽ)^�ȷ!�T�д���\;~���ء�Rr���?���ؐ��d��!��&���r�Tc	TS��V�(ڲo�yq���?s��x��/L�%1lڣ��uto?�	�NDՆ�W��Q̟ܞ���;����;���Wb2���e�}
������
�A"�gJ�N��\��S�;�Mk#,�ȼ�sb:O��@S��ѝ�;*6��U�¦z�`�����^�;~��k ��ۇ���sp�8����{��F��Q���E%�T��խ9�5tB�RS�Ă���\P'�Q[�yI�r��=iS�Y=Â�\[�<}��]h�҇�t���Ba��C�Z��l~��4��xg�%���������~q.�˃�@�g�H���|���f|����݉�:���CL0>�w�$�E1���;���E1�_?`	����,�iPs0�7��6�K5��/�Px�n���T	sM�۵y�|.�y�7�M-�I艭B��=[���"7�����`�ҰW�y���h�%p�R�,? �7�ַ��\�]@\Hs��c/gM0m��?;%�ui��\��A�
ĸW�����XԖrlf�P9�Y ��,�Y4�u�6|ppѠ64�ߟ��\�e%�B�rX������9�b�.M#`��*����:�1!�r&ܧ>y.=g$0ǝg�=Max�ڞ�c���Y�=)+�6��=2�Ĭ���6ɤ���kpL��4@ާ2D��#䏙���|~����ꊬ���s�OcV�B��-a(�d���m���T�?�w�*���W����3�����t����P�����ɣh ��}&���aќe;�3F��g�/I�jo�0��y�D�#v�\L.+?�0��v0`����8(�`G/�]Q���R���ܪ	�R�����E@��EBJ�HE�h�W߉Wqt��ۉw@Bo��o,⃛ɼ��]��uTY������A���:3nw�Y�(=�7h�}і
x�Z�b�K�ܻ���ܣx�36o�R�lcS(J�� �̛����o��"��x�6a(z(]�Q�������,�D�ڰXo�}��x���"_yJeD���ڵN���
��Kn�BfgN��!�/�s��1�f�!4w��C|������0���~�7;u�.`4���
�(�i�Y=o]���ծ*m��'F{q��?�Y���W�9��P��ׄ�g�`QTs�)�(�\0O��@�
r��>M�G/	4��"	w����E�7)��+�|��iQ>}u�
���Tt:`��P��w�C�.Ywu�&]䚡޽���FO~X�N�Ȁf���	#í� � �~x��T��#j�=�����K}3M*�Zd��?�X��܏`Ν���b8X�l����E�駰�R�rE6�ߣ���X'u`�X����
��l�,��r�	�Y��`��T��ha��Ce����� =�����̻!C�`��4����	&οrt�E����e� �������ZJ�#u��S��_�#]�@�T�l���|n%�����r�נ�u�)�X��
"�1-a�϶��u���a_��	R� i�j�ƩMod�����̆ղ7L��wl����A���6�ԃ�v��6���� ����AF�w]�u0T*�oz�%�_��6�;T����nFt�Vl~E�\�
�Bٽc�G]0��� ����V�Q��N�e�38>�^�w�������7��{i��i���C#C�Wb����e)Q�q�?���� ˃ݖ���N ���ea��~�a?a���%��L�����^B[?������=���LsbZ�~0��	>A�<���p��(E,�������J�����,�UY5h�ߖ���r �����i�]f&^�ڴ�4���S(a�ޭ*#G�8���Li0(+�s�æt�Z-(�W���./1�� L�Dn�V̈9yQRf�p�o�9gW���RR3���$�N��QT�N^��M�r۱��i��Z��R��b3.�s-A�W��ڳI�=�c���UL�Gg;�R�za��~�yVth�7Q��7}���k`M���{��҃�j���C�| !��p��o���g=|�����]%Qh����A����A�3���j�}���!�/�I�2�ܵ ��T�b����S� �
��m��ܙ\&Żs��((Ɔ?�b;���[Abkhߋ���i5�4]$u�M&��v�)����6	HI/���S�<�X�ޕxZ������y��G��j���O8����{͇joG����)�>,Ly.���"~p��]����jB�S^����d"g��`;�dBBb�?(��!����f2a���a��s�$7�x����i��Z���OP��,���|,|^~<�A���Rͥ��jh�M?�͢�R���{I�j8�������y�g�̏��\��Wf��H�o6Xj��/p��ܟ�[��2'��y��8.`�d�p�u�0����M�Nh���B1v�*��/?&��,�(&WD>�rT�v�E��L�9O$��*l����ɾq/��`�0@�6f�_rD�f��f'�n��5�(��B$�qcb�5o+��u.�(2��vv��-��s��|y~}��H�tO~��cHHC���1��Cc�C�9� O����PQgCa�T�5lP#�z-��@G�����E�4_x;�wv�j3Be�c�7�!����O.��׾�n��v�xUq��l�۩�S5�,=ƹŸ@ g:67�!p]v���YP�6�a��)F~�C}3{J ��R89R#>o� /G����[$(�����X��c�8���,B�T2^^�!��A�,�ؙ�T�0�SE.�|���t��h�R;��A�Z�p��`��@��x@+&��b��g�a�)��1x��b)C.������1�<E��jY5N�^
����ШT�$id�14Դ��=�[����F&|�j}h��<���̚8`SV��M"���x�#ӌ3°Y�I�NmvI��#m�V}4�|������	�/%��Z��D̃��1V�~�����
�5���_{ܾ���Sm�ty���	w�ȑ
���'���+���Ō��&乩��� \�ꝰ,9;��no�����U4s׎ߐh��N�E����f; r��1�R?l%L��>J%."��bM�TCLwE�ڗ�j��U�E����1���P>�S�|a���0c�N�E	#�ۏd��;����2��*tu�|�V�+���"ڃ�r:0��A]�&�8�A�^�5��hC ���/� �	:Ȣ�o?g�i�:�9�Oi��nBl�r��Ġ��p+��c;i`GŰ�|1;�bq��9W�Զ��ȦJ��ɳ*Z����+<���[�����}q2nl8����|���xNgq4\2*��]q��>(#��������:B���\n����<�J:�J����>�Q��|b��n�r�l)�Ofn��x�>�@��u��\����E�β�E�@050|%�i��;q	e6O�3�;�a�5u7&,v��$g+Z���"bnӽR:���;.����K��t�4��_���D�#�����ᘔ1S&�E��c����,oq��ͅ�k/J�.��K1����²��vi������̈́�����zr��>�;1��R�����͡~s�YQ�jN, ��m�fInҫ��l[IJ��6�x蒖u��W�/
�ߥ���'�K֭��=���1����:j����D�J
��T����l�Z>��]1א[��h�>A"^�	̪�O�	����\ع��D��D��?���.թ�����B��2B�;��9�kZ��Pʹ�'��/ͬ��9 �{n�K�Cӂ��T����zD����,Ŋ��*��UO��t�9�=~A��`�g!�N(1v֗��_˯�\[���u��������� (��j�dX���
j���R��m�C�w?�X(�K����B�D(6����̷�=L&k#���$�ٲͱhW��_�V-�9j ��u�g��B�k�%��z*X!�}?	�k �C��^��߾vM�h�qc�j|ݺ),,,���b�LdtQL'a���&��,�����C��~�u�G�Z ��Ɂ8�B��� ��k���HXyxR��-���%r��mQ��v(�+.��R\�
��T~��u�E�~2�����	��K,/� ��弒��;����V����;s>j�X�
z��8>�%@��v/��#]�*�_��XD����Q4�ٺ����L�C���I6w����Kl��P����\�ޛ*Ɠ�O }��$�T:���L�6�K�����ǀ;��G��r����*cb���=sF*�7�d���VP�F�Q����YR"a�S��󒈿]
�R���z���[�]�`x����ٺ\�=mL�b$s_c��;2z�<����f,���Z���J7 �ׄӷB�/u�Ҙ������W���f=�P�˄�6A|K��C�N�����T�$G���mA_t�m!��5�n�a�7���ӉZ�E�Ü�9O[�`��X�4t_����h��ާ[r�AaG'��hޝ��˞z2g��*y���c�:�Q�����oT����2�f�h%�A<�n<x"��[J�����A��$��!��]-,�h�jV"�Ɇt�\��)������!>g��~��ƙDv��ى]�Pz(1���7�<}_��9��I� )�3�6�
�Ǣ�t���7�������(��2UO������y�?C9�@/
���Rx�߳������n1uY��Z�(�R;`N=�Aa�Y(e��/���HN"d��a֕��Q\��Z����W����B-��B��8%R��ޥݬ`��b+�x"��d�(�	;G��D̐�C��]W��$��+���6�r%�md��-Xxg����Χ�r����� ^��>��nСcg�o:��� [������2��m5LSD����'&:��h]3�^�dt���Zzc��]_5��b3tc:\�#�C(���Vib\d����{]���t�P�����V@z
��b���>����m��[�3P�&��;�e?�e��>� �_o�l�����Jj�ƻj����.���'�|�ʇpHX��?'o,'-DU����]�����!K�J���9W^�F'wF�o���,����xVPA���C����s�E_�Dh�f�Pv�����Z����j9��p�j��G�*��FBfb��N,�Y�6Rgb!�����Q5�,�[e|��*�cb���%�2��}�w��T�ҡ��N��ǘ�vЪ�ZY(���{�ߡ�����(�LO�������L�,��ï#Z����(���t�O߶�'��/˖��4����B�f����
ڜ�E������t�qw���g,b�[�4-Z�@>&r����Ub��d��_������8���K�H^&���q�=;�dw�8÷D��B��8���}��;�T��K�[@�5�<��O�$���j�؂�[�Ep�~W>����vdq5"���욾�����U��P)0o�ө�ӳ���Ͻ[��Î(�I.D��x;B�L���ǥ@d��~.�g�J�����g�y�`����%�RN��f�Qw���e֋�D����o'�6�_OQ/�RO���R����~����R�x_h��� '�q���T;t��nm�
���x�p,�.}��!+���P�a�,��#�V�G[���d�b�bL0r�C�)8�g���t����~HV_�C�n>O��=ɩO���Cb�$�����z F鶁xpX����C�)������6�zm<�����m����Ŕ������� ��S}f��fe5��-��ezr�wA��|�رY*� �d��E���n�\�06����(]�o�J��z*�2]J�I�)�b��Y��G\��&������:�x�7/\Pn�bx�W�Cۙ�Z'���RQ�BeR7����D�_��Z��坕����#�2ۊ�`�����>�E�Vߎ�
`ME{�5L��)��h�wI���@HA���i\�J;�w�T�9����-o�"} ���_�\�jo�Q��V��х�30#D�0���̞�����x��u�)hz�Dh^a[E�\sǓX��w�d�n�K�l�d;M���r�/�0�#H���4���>i���3��������X�~�M�Òr�
��$u+`Ҫc�!�<���&�9!���Ɉ�J�!/�6F6�̱o2��d-���X�+]K�P��)�!��U@�����n�P6�?_�Q�����z�S��`Y4�Jvn�t  |d��d����Uo�?�l_�&f��k��_W�w��Y/�@�c�nc�^��i#{����R��7z�ж7�N,�g.\MU\Y}����&O�:�$���PIX�G���z�X"����6Rb3X���l;��C��ATv�o�P�ب���>���T��O�Q��A]L�[}I���`���T�⡩��D<''At���*���'5Q#�`��
@Is�0��R�}sM�n<��;_:e�lT��ʸRMo]���ŉD�9�/�M�t��ðZ��U�2��D{Tp���q;@=�	R�����]�K�ʺ�6�E"������H�n�"8(Kp55m|{JIb>����T.��76*/����;������C�nj7��ѐ�(�(���Wٷ��d�ٮ��u�Y�xٽ��'~�tJ�.��&��{�G��d%�=�����Ae��R�_���sś ��\~��G`�e_y5�I�2+���8�{�F#�c�ƲQc�P5=[-��	~.�g"�0�3x���%i�T@?�-gi}�Z�i�C�>a�('�|J����,�Ȑ+=
.�gęy,�O�K5��:N��j-���nӴ5�@���>K
��0�"ɂ��ra�ʧ^�7V"˫��w�@�[WH�@*��p�Bm�Y�!�y&�#bzX~��[!�iy}6 �L�6�GAN>���K�Zl�DK����gD.t� K����x�gO�y#p���|���w��QC��E��ϞV}]��fB�u>+�ٷ/���L��s���=k��L�}���i��<^DN��J=i1�/-���؍����b��MW-�X��P�
Npm�(M���A���!�&�t颲9R��#�'��OC\��#w%��[]YȘٻ襯���J*Wy_�@d_x</ຈ`%{ �C�s��B��������h����e`�e�D�:Cp�˘j�*{���7?M�m$d�X_ �3$��?��fd���T�O�HZ"���t�B�>v�'�3��5��f�R� �rn���T��Х�A ��ǤI��J�pCNn�ʄ)b�K�6�ڸ��%.�v�t�G�ZX[sݯ;*�ęU����ɟ7)��ܭ��J��+�/|���j��#����i�.d�DFf�8�T�֗�4-J>R}ˋ����I[�cΖ�yu�J�6����B^apBC�ʍx^��+�1Zo7�t�8���D�J3З$t]���i= !�ig�>�';�ᜩ��� rʕ����c�A�q��K�o���͈�kq�Lf����=���K_韖E�{��6a�%�?}��R��?Ǽm�5<��mv2��Z��}���Dig1�)Ά�4�H�=�zw�Q�#��<U�[_�W��B���sO���@�Ǧ���G2G�\]2�VL^s�VV������{�I%��_s=�o��:y�6�!�9�r�W�(���:]1�s�[�C����b�/R�������︚p�8��ޱ��R2��s��XƼ�����?\Us�2A##�^6~��bp�+B�9Z2ݰ����_� e���/i/�¿UP� �O�ԛ5�"`��'�`�|4/���1��-_B��ü%M�Sqv�'�)y�M~��#�k���w8�����-���T�����U*n�j�daQyhS�Q�e���p�hΚk6Boebٯ�Ȩ\ԍHp��Ӑ��w���>�	���3����|����F|c�\����l�è��\��q3��O�â#�\�a~-|NˋJ����Z�>�^l��`X*���;����爱l՗���R���s��= ��ȯ .]���w��C�Ux�M�� ���Tѧ�E���O� "����5e��j;	b�/&3������,GΦ0��WP$y�.}�V0��:I�Fȵ`�V���)�7v|� �Q��Q����н���B�`�5��r�s~�n�l�!G��O�:/�=T�N{bP��sY�����1�3>{~��̷)
	�'4��~$����l�U���~�v#�,_���N��.�\��Gǁ��5",���Єl���eW�l��G�&u��N<�<z�PS�݇`5(.|�S��o�6j{�h5B��T�5��i]xq�P#���|�?Cs��&�Ns����� ,�d����_������/�U�:��v�稷�7�n��0�Ɠ*�7+����0��K������*�t]@ձ}ߦ��3��Am9���7|p�	Y�����u>.
g�<�z�Te`��zJ�� hd��_le�2�:h��+`8��L�?���Y����j\��>b{���mH�]QBa /���ڼ����"2��o=^,Vj�V�66Hm�V},���NTt�䉒m��"�73��54��`w�`f�kc�_E���_�+���l�R�O`H^��z����%Q�
�6�z?IQ����r�kb��|p����H��rs�+^�y��%E~^%r��,������"�<�n8��$m �hՙ*���g;���Dq�8���.3\����I꽎�ʂ�c��<�Hg��iV#��/<�E�r�*G`��:r�:����>�+M\O��}'�(�0��ϰ��}M�#������~mЇ#�h6nJ$�)i<X�ȹK� :���\���-)�� qW1`�ߘC¸Z�y�c�Y���7�A��k�1�&r}�v_9y ��-ƽd��B�����k����-`�e�o]h��)��
`��ͭ�](������4�,�d�~:E�-0F6���'4�_��"h�KF�O�ITcWfItG���
�HY��J�3٦���'�K��Ηjd=���?�|R��TO-��)�����w�a~r���#������6	��%��#3%-*�P��l�ۓ���ظmq�M�1]tD�4 ���>r1OLE���@�	b>���u}w�G)Xp�����	���~��/:z�ah0x��%�����ѧ[��{C�����GL��7D�5�Hr��B��WY�YE��xm3=�~:q�"�G�Y玐�s���q��`����c7��|0閒���!_H�P-I2z��=��Fo��t�]�x��%xd�Oxv?z��\|�ψj<�e{��n���ۺpw�Sj��af�B�[�/k��f�E���0��vj봶E�|�Fv�Nurs�+�.k��'��S�	(�` ��+�ړ<��@�|Z^í(�l�+������6�dh�͖�����AN_�A��~�1�{�[�7�
l�����b�K=�A<,��>S;J�L�p8I����9 p�h�̮��*e>�������˘3����bv�65w�wj�{���Z�m�֛o��G����/�� ����l׶G:S� �����4��5��{�[Z����n%���Z���POI&JI�G�ǧX۸Li��OzM�M��I�:zPAX
�}��o��?E�{|�/j�U��k�K\1���3������l�P�M��L4��b���Ԡ�ͤx9żN
Ge4�˶��m'l�3��{����4���O�旰H�x�
n�ӛ��͎��Қ�2y�7�ٕl�djpp;�- 0��/����k#E�I+���R�;&��U2\��.�a�ۺF:��5����x`��	��i����r�"g�{�O/u�ι�!T�3M�@���/ύ�D��n���uJg�Y�r$��>�+`qF���3<�� ���V����T��oż��/�z�/�?<�]&ގ�$տ�	u2����;��F&�~u����vf����}�0�����d�H�_���'�N]�EU�|�{�W�<�&�q?.�6������]�k�[��!c~�i�7��Io(����|߳;��s�^�S=۠���:
��w'@i����+e>��������-I�I��0�.]hVNM}^���Z	�~^̸��;#���{��V3)�SHmk	��1���*q�u� d͆�9.p�����,W���� �Bh/�el���&V_��,0���P��"�f(.>*b1�Z�ž�"i�r�����J�V����ſ��m�@�܍�*G%���u?-��k������rf�99V�7��J+zBh�3�Yd��&�����C�f�vU�"��<������Y{!�O�7����gha�f�[^3Z_��
�-txr؜�4�ä1�/��	6YU�Y�����FlaC���F��Y9����4w'�L������m_S|���t��j[��\!��3g�P�����,�/M�a͙.�y�$�q$�YS�[����r"�zv�՗�[���� �A���T����R�>��V���O���p��o|n��O-�������>�S���HN}�J+���5i��� �c�i�}�
g;�z��K5f��aۯeO	���}��pEz*���E�aw=�v�b<ϼ�b�3�O�8s�r'3�j싶r�6<�u%���?�~�U4��)���&R�����}%
�3CW���sC�8��<��	"�O��B�>"��9Rru�3�v�/�|@�8��H#9�y(t��$�	�~Ŗ�L��QD�e�\M�tr���@�d�0ޥs-)޻K�Y�����R/�<j�ξuO��xc��(.�㽪���:�N�ZP�;��9;����BC��Sp�紷ʖ�<���u��)�-��YD�c4ʦd�8L�.��.�u�L�l�F��1�O?���D��*��C�'�b��w`fH���X���=�D��U^���Q������1y�Rmpjw'��z5Ȟ���O�!��P�9ZH�`0�ѱj��5�3���2:�)��r�Ǹ����q�,� ��{L-V��w�
������6jb���ΐDWL���X\7'\Y%��QDa6 ��3.,�9�lP�#�*��g�ߙ����1>�����p�娦�p^����A^��y/��Q!�������=�T��K���8�+�*H��'�n�(��M
i	,A*�@^I�o�\�`I�� ѽk@�K���-;R#���F0�z��W'TCH�VI�x+��� k�Zp�ڙݔ�DS�Q�HX��6�&!6^~��\bq��t��x���������7��ѵV-�>��@b�ì���t��w��,.@㉣Hb���uVo�w�܁B��m��1��j���bkbk�m�v�猥+���W��h�{wѧ��7�i>�R7aHNK�	H~s ���V|Hj��m�k��-,�l8k�Y�Z� �6Жu�Z$h��Ta�ٝg7'�o�К��J�0����\���$Hln��}���y_v�>WΨ&�������<=X���m,bx�.��H��\���	�<���3����Q%e�[Dmw���~���M*w*q;�$!Ī�����,�և�`܇�|y+�*�;o�%ƣ7#�F�|:4�n���pJ�T��Kn��� 	6b�=X�	OH�to�9��X���7�(E<����鳕�ه8T��4�G+��{�%�exX���mYU�V��:(|�����"�lD3��H�͂�������3_,Ŋ&r&���N�HfF"�#�Uò;������9#�[��B-Z�1��"i~Nܗ��'YO�>��f��w�ޤ)�w�E(.DU��A}ɑ���f��J<;!A��n��rsX��&'q%n�.��s�|�"ƺY�v)4\r���0�bĚ&v�5`����֤J��:��� ���_F<�ѻl����$��9��g���>*�ͼ��� 1|����Y`���奢iF��n�����f��-�z�Q�k���[H�Zȝ��f�\�e3�*7$&����G>��]��e2xJ/�ZQ��=��)m�K!f`4y���B���~�������_�7'/L[��ErR�$G����~Z	�a{J�o߅o�8kJ_��������2�l�o��鄼4�P�0�܀e)���vȓ�VK;��ܽa�RĿ��儨e��,���a<�.��p�E��y�,Pj�(Ch�˃�)2P'ƍ&�A�g?�h#��}�]&!8��|�=:} ������k��2�-y�"�y,�y���NqJ_��f� |���#Ģ����IRM�-&n��]��<m\n�򘊟�\��z^��\ᥰt?,��d�2�6�>F�K
B�9˅mDBS����@vE��B��Ç�!7�
�ȁku���G�Z2
ュ�(����-8��a�o�[A��i���eW��$�-( :^���	�2���Hg� "$9������W�(`�ȼ�¤��@y�M܉ȡm����"#�M��+%n*�=��biX<bcw���^�^���O�T	��灑��oG�b7�m���1�Q�U�JQ�{$���ў��lZ͵o܇����M�{߅/��$�zuc,�uS_ib1�V|G��F:�uf�?9�1i�A�*�5�Vw �;�1���k, ��q� HR�0&��7?ç3C�Uc��e�p�%/���YF%T7���&4K�Sa@m��9W�1� ���j��QS�A2���ņ�B��jw!������P�9� ���aw ��@�SN<3YI�=�e�>+A�D��#E�������9����}�v�d����[�T�N���r٩8�Sc�H����P,ց�s�Vk�w��,�\Wn��l��R�� �5�7bpս���	+�E�Ev����/�Z0Y�q�P�Z0/��`�b<ӡ�Z:��t��|��4�`|�e5�1�-q#�,���f[9}2����6g3��0 Y�K�G�߶L/�n}��;N�c�r���y9֡����F�0GSf����÷�y���Cjmum�����:G1_|����^{��P"��(�[�!�a�th�o!�VJ41K�3�1�F)�S\�${'���T򗅢OM�<&�&�Nj�Uk���+?. D��>��V=N�Q��I�E�g��~h�
uGM�.�����VZk�R��c�nA��r=����3(M{H��Ngth��5��ㇺ1�_����`�.G���4����1ﳜh"&�%�]>���CRW68�lw�����9�ja�[�ey�o��D��w�B����%�Q�cp\F��o-��/��)�EU��0i+�<������L$�v��<+��1��x��H>�x��c����agH��G�B��~|JpDڙ̋0��Y��;g�΂4���de�˦�f3�������#m���w4��#EEL�VcJ�ȝ��=��@���O'�s.䐪��e5�T�q�D?��b&�a�SbaFu �W���U_B���[o7Z�T�e8���e$��2l�X��Y9���o8y�Nk��5t��@��4ǵs�����~VzV�s*1oȃ*%���g���i�U�S �d�\ۭ���H酯ϯ�_?1���O�� o�����;n&2��u(���;k$���*�Ay��K�Ga�& 5$|t��
���K.�#d�ȍ�m"/}�����aS��h�&���^ֆ(U�����Dú$#Z������sP�)֙���#,Zc�\���+j��g�D���Tw��	g(/�5�� ��0rw}L_[�e��ɟ��/��02%�� �1JmW�� "p�o����Tj�M^��r�)�&����u(�~I;����� ��&���B7Ґ����y_���Wp��t��#-5g��t�P-, 0���'kO�#z��&����s!�v�h�6�'+]�"���_�ZZb����ez�.��ec�z��ve))|(Yy����5��ߘ`R3Nҩ�V�ַ\q��^�1l�TX�o�Ri��l`��~��S`�����μ$�K{�;RE+��Cz这�|?�і%k�l;�2Ù=��ϫ;��%���ڬ�屡/�,��|s�3m'SZ⿭��f���;���R����BɌ����T��@F���Ǩ�G�O �+�̈�llw�,��B��pU���A|���~�*?�C��LL2UͽF��ñ�G�.��E�@@���.�`Q�?}G�}���cD��a���>SC���( �w�_Ѫ���G�hՓ4p���t+���n?}EM �d�C��93��<j�x
�x&8ś���;:2��w��ԛ+?ڋ��K{�r&-��칤5�.�+2P�S���_ְ/�ߎ�Vƫf� >-s]|LSV�=���֨mz�*�$I�4��5fa������/_�Ϗ�h���_�#~��T����}���BMxT!p�VƮD_z�����'�0��4�/WLi����k��C���ٿ_/�3�_�:��[�7�0�R�v����ђQ����C<b��+��|)����f0�#6�_~fď���?+��)l�)bkO�ըX{^6<t�W&tϐ��@�a�9�(Ajm'�t)
��J�S��z��`mڧ��$K�F���g���A��҅Q����O�-8	pK6�bF�P�{Ck���/6�jz�M5� �&X�)7���#��-�֚F�0���:��*�g#�;����B��5uI�4-��;!m�a>�&~W���˳d�o8S�c�~[r,nfM�p�����5+J��:ܸ��P)0�`-CL�CX��=`�⿌:<[�����)��S�"�ɂcRs5v,���O���#٣�NC4��mC�3��8��X;u��ɤ��Z�W��Wd/���
e�Qɥ�b�8�ݻK�x�ܷ'��D�;�U�Kv�{@��>7�{�Z�*n�>(��ԶO�/��7!�6����@����Ay ^�� �;Υ�1���Ӷ�P\Vw	�����H�A��#�	Z!\�����BV<��:�d������j7���Yi��O8��3l�ux��f���-�k)�2�Y�E��.������}3�=%���k���)Wʤ�29$��u��E׻�m r!��<�:v�ٙe3vm
�K����h�z<��,�}�X�jADpG��%t���<~*f�[�̻����� ��$6X�����
�Bzg�e���7�%���}L� ;�Hf���1�ӏ�t��G~{D�%6u䮖��D���+��q�BTz�4O���$���g�!r��,v�N��4gb�r���eB[G�3W��O�/~�Ɣ[}�-]bI49��X$R�R5�K�O{�P�Bx�w�1� ��e%[}��=w��R]Yg���x�2s�^)�Mi�*87+�(X~�:�S�GkH�RfM�𺖴�n��^N~�g���O��Ynݓ��ʑ(�����X���h)�=����W���D���șg�h���F'Y���4���B^��������U�
��US՘�_ ,^Aꆀhu��p7M�Z����� ���{w�~K��rτ�K "tA����ߤ���P`��͑���	#2�$W��r@5�9j��Ѭ���JHbzk]�&�l,�³��q�-�u��wh&��s\$�A q��S��?��lY��2�c֗r��p���܃�m�^����X�=`ףT���<H��ه/�����[�>��6�y��9CK%E~�>5�ln#��N�_іLhb&v�w<�=@U��oJ��H�����Thc��<�Q۹�+��|$��v�ʔ
!�8������	�
dl����Jӌ0�Ux0��j�+�����+wy��k�}�{�DK7�'
5Ere��U����(2<e)�h�y�xk�T�<`FD@n\��7-�0i�;�o�~;n*	3k�#N��߆�V�f�-|�����9
���4��7!�q�C�!��vrws>����������5C?G����}Pa�I̋f�,y��*�Jϛ�A�PFN:�U�̯�`�_a!(K髧��^+eӽ��D޶���
��|�Kw�/��m�R=��	}�xvL���U�Bo44�Y#"�ך3�\7Zȥ�c���]%�X���@ƾ���(��)���Swi#b��v�����3�W����\��"�����)�1^��þ8���b@G$[���z�O}���b18�,��985F���H�;�Ғ�{~��։�a��V&Sf9"T�NEC�'�W={�������4wWp�~��N�C�C����`:ᡬ/��LȐ_�:�OPP�2w�_�o��xG8R �ފe8"�'7�A%�!!���cG�@K�Q]c�1H�z���u<�ai�?,���2�Yh��ي����e/��)�|�1WD6)`G�p�k�����GSDk�ؘs�0އk-�PTΤ�1^���q�Xn�b���puGj<$& �tN]K���Rr\'pE�r��e�&����/=� �[L����h���7zJ�#��*�<�nN�|�s���G�^���.m7�5���{��~锖D~6���H7Kz��x鐳���;V��Ƙ���ݾ�������'����OZ@yj�rrs�?���;�|C4`&`�l�R_��C�	sr�y"�m�Q
xij�1��������F���N�/�.��lF	�^PՎ�DKX�m���l��<�I����Y�"�_��0��P��@�a���g��V���Jd���V^�*A���D�?�m���\�6,�5�nw���.�]>4�EZ�;�x���,T#y�S�>/��3�:�����@3�^
���"X��c���	�r	FYil0��$K^���l�_f&F/T���ڨ�)Oe�:�e�s��l�i��{i��b������3�f�4 ��B� �����'�)-Dٖ�R8���7�L�����ƶ���?����>O5�`�	Ne�{�@T` �XK�~2`�١�y"I����Ʃ�����h�q�i>���h19��kB�qp�/�	%7<����h)5��+6a/�e�cr\FZ�R�'�d�5s=Pe��7�<y�^��wxA}{��~o!oS��3W��L�E28O{����gZ�/�_�:v�n^�Qn�r����Qc6o]����D�q�To�=��]�	���6щ���a�"���YC~�ߍ~}kL_hϯ������NJ��w^���^W�� �02�7�p*�(���n=����mMe&��u�3����t��$i�Ԧ/��z,3��4�7������T���F�M�GB}7�?�}���6��<z�T���]�{<����4ܯpsSr������S/F���K[��g-é���7�H�L�҆Pv�Ce��,�ND�޼MR�ȹ��-�ğ�R�Гv�&t�Ķ�2τI�w��B.��uf�2�9�xFQq�ޔ}L���&jK�]0���k��=��r�`�BO����Y�K�$���<�L�&�Y�̀;u3�>�,�U8%j�1����p&�hk�[C�d�Dd})Ι�>Y�� 2W��SG��9��C򬁉9���Ts�������~]'ԿB���Q�TBŸ{�U�[J������!R���1�����D���ɬۺBF�!��������Cq��(�w,|�@�4�Q^� f�A%���ԑ�8�<��x^�~j�Dd�h�TK:Ŀ���.�)z�L��^���19<^P�5?�k�\ha��Q�ƉF�{�Qq�	���� �e���@AU�.�ϒ��b��n�-bP���Aô( s����2��50r6h�l�����3X�$Fu��$�m}���ѡҵˍ̥-⫚��SЋ�J>nL���ΆȮ��Gh[F�<���`�[�[�vDꌔ��4P8&=zU�d�_��o�;Ԋ�s	$vRT��2B���4h�����2<�i�&�ZH����~�o[�'�Fg�Aͻ(s=I���HUʚ�R��l��įmʐ.[�h�����J���i�U���ZK��ɚ|�2 ��>�G�"`'~� �#�ֵ���5�ɢ�6q�G�(& �F��a��=2Aq�6�h�j;����t����l�A3�U�V.-.q?Y��:�oR���ڢyc��:��>�c���ޝ�/�&T�
�=����U��B�~�ݳ�,c�Od�s��*�>�Nb
�AGꈤ@\��.$7�v�t�j�����$��O~����,ǳ/�)�Qg��Wm6����:�T����z�&髎p����B�>���"r�dh��%���]l�ja�S�փ�8��5v*z�a��,�;�3��u�ms��!�e��dm����r���
:嶢�Q��ٸݳ���ܗV�/!0;���[��O�!�����߭M��=گ3I3~��\�R�ؓ�~�����jc+�-Xk Jr]H��O�������i$>R�	�tB��vr4l\�zN������L��f�r����`���i�"�r��zJ�u��;����:�?t
 y�;r!�/���6�5�߶Yb�0F�C���w `�76w;"�NGݖi9\��Mf�:�ۆ�Iz��u�	��"1����"���C�j�$�h������������Ĺ�^l[���;u���y#K�����k�f����g'�y"��m�D>o��4b�����6���yetF�y����dp�f���-�H	�[�� �N����!��{RJA�Y�G�~����������M�OZSRfD�e0$�>��;ׇ��'��J��a~
�`��z�l�c�"7ê�O�p�X1�Lw�y��3NSO>܏4jt��^*r��¦�X^Ǩ�a�"������U���D��+^O{��޵���8~ �ޙKVS� ���O���˖]�wHe��j�Y6�n�Lb�N�0τ\��:���0�������@P*B�3���iv �3�N���+���	�����ER֕�o��w������ֳ�|b�P�[��a���=xޘ�w�q��˱�W��[�s��%<��\��Y�¤v��}.�h�T�!��l{!�&��ʘ�h���4��2�v�����1S�Q~��T�9d�<���v��V�G8���Gٔ�v�^i��Fir�yǆ$����/z".�Q�UX���0 ���d�F�9��[�M�p��U~�C�f�"}�^w��8$�Fq$[�VFB�+Q�q��AA���tz	�"�%�h��4,�ҎeVc]hJ��)e��j��z9[;&��ʭ���r��Y?8m#i.Ձv�Q$�[�&���LX0�Za(����\��'�c�y�ls�war��F��oo`��y��"��$?�P"�Jsݎ�Q`R���̵�)ʬ�+�F�y�L��_�Yc����g�7�o�U�H��ߴ�9bUR&d+`>�3�Ln�h7y���������lQ�r����	~m�>Č5K���a1 ���i��܇?c��mjS߽K��܅�4�@*�_K.�z(�
����ɱ�7:76��S�u� s��Az�:�N�C#����$�$N��>�-/�[�2o`}�W�����2r��C#<笖��.Dn5:��<2�A��
���A]����,�3̑�o��Jԃ�(-������އI��N�x����i�j�����/s/�͟/VG4�@Vf�4�z��|k�5�O쮑ö�Hh	:)@��Z� ��0H�n!7�������ئ�����$�{~�I�w��f��/;���_�P@l�Dn#y.�;j��\(���������,c���o1uk�b�!C�f&�X_р��D���G��Q®Јp���_�[��X�<"�G�A������u����%�>h(�D
��}�uk�}�h��I�����S �u�|��IY6����.wi]�YFa�@k�X���O�h4r�8��S��R��#Q%���q,>����7��S�E▎Ɉ3�,�J��Z��b����n��TB���p�!Q�SF��æ�Y��{r7!R0��Y��x����jÖ������離|��;6"�/D��Jƻۿ�]`�����9�'��գ��:7��6��V��v7�PߵgU;'�¬8�+�pܛ@�\�I�dV�b����g;�9�e�f�)��'{�1\-�JsD$]QsU�#�d��"3�	|��,ҁ� exT���~�=)��˲�NZ����;Uί%�����}�$7������?�zAd���X`E����&ּ]�e�R�;o*E?���d\�3�"\���a)��K�$��
!�K��=R�	A�pZB cBq3{?qm���!b"
�}�u������������gsX���^>[ ۟FH�?��Q���gW6���YY#~�	U�~q}~i>�]� ��,�d�h;t����U\����i|����&��[x���Ø�-�����OH��1n=����l{�hI[��S�)I�����N��K���O~2Vsm�}�4�Y?�P�����٧=|�rv�A�8�s�-M���w<"�oCb�*�޿Ҫ؋"O�m�P�oZj�+R�0
���&&<��Z̥�~�@~�i�fzĨ�����F7s
�e`*��U/�g$��B(ۤAXI�H�~�l�%LQ=a�$/���팥C��U��b�,Wݭ歆(��ȴOc�^b��m����3(��R������M杙���T}������x����sg�H�+����ݟ̖&�'�����8N�Lzp�wo�×?���R����Ӻ {$u�A�f���0:� �Dq�S�U�pI������K>��]��wLWXlK�5G"@-��Cœ?�[�&h6�܇�@�$��
��a,����}9���#�3%��w�������0E��^�W��;j?��؟%K0�� %���0�H���2��e� g�g��;�#,��6���P�o�7B-:
VF
�؊Ά[�G�Y�[CbN3���]���d~L�o}!�39e��S����1i�8p�)���?W�Ɍ&�Mr�E�=�%��������GO&^�K8�wҟAAb��9�"e��#b߉�d����l�{IN�nHw{k����Ex8�ID@��M��Tn���

L��LRS?rA��[��ҎSq�+�?�9�+U/��]F0ˣ����=�;�:�u3%��>}�T�n�ڵ��!�hY7s<�_���/�6�^�?m���U��>)��_q�w�
�ZLS2�cD��z�T݁P�`�-S4�D�J�"�4C�q\�]��j�xN�ؔ��� ���J�(E�S�,�ݟN�4\�F����{��]��uk<��rƉ�v,3Z�8�{���T�9π��qr>�
��$	� �-��y.ԨU��A<���m��������N`��Y��׺j�)է1|�$ ~@ŴG��qɨ:ES�3�,����Z�+C���S�:J�����U����@���#	���� ������U�1��$;�G���'�/Ztq ��}�'B�^h��^��}oP��`�46�c�����k�wq��W4�lF�؈����.�B�ݗ�rƎ:�.��.K 1�
[
�?�;�U<�P4�o�d����[R�����V8��-+��O�
k˞#��Tr�`Ve
>�0��|Z�������K��pN�1�� ;���(M;��q�x/��*���{L����mȊ�9`v[ �p��#��cIn����n͇�7�͹���A�>��U�I2�L�ퟋ���m��6.�{����f	�l��s�*%�AJGf"���?/�����S�n�<��y��V
�[_IF�T�s�w�I��6��z�Hc�\���^�3rL�*�EM߇�T��4{jK4�
j�/��/Ԏo}�lG{6m��`r�A��+��ce��5RM|ؔ�$e�vR��n�<���[UZ�~��t'R���ic��%n0vmK���V;t:���M_%���a�����DF;��R�q'�ү�;��3d>СWI1'?��aXݙ��j�#��]lmJ���V �8�m��WO$/̧PR%© �oW3�w�o\����3��������˪��[����e�x�軪q�z��XP�l�AYAHA�1f�ࡺ[��_��ч�ie�֥[�i�k�Iw��26�������|D-\%-(�>O	2�헇۔E͸�Ln�ɲЖM7��b�t��$�W������F���=�}~��:v�Du�xs͞2Si��Mr�q+)5��?��h�+�#�æD[~�����qo�_��>��4�e} �e
�/�uF�Y�F���J��fF`��wً��zF�|��D�M�ӫ�j
P�6�P̴��ƶ������p��A��n4w�yϓ	=?��� ~��$�AJ�;�DX����|X�"|���jwPxA�أA�.m1tN�y�ȯ{1���Q�	�H"����[5^t/K��I�齗��0S����N?���f#D�d��q����kv�X�g��7�G��lƣ�9D�X�6Y�,ge��h8G1�@�o�v�G'�a�]zy�* Z�b^c����U�$(�kR5kF� 9U;�u�y��k�B4���ց��0�\J�z����n�	�Hqٝ�lr4*|a�@��Xf7�{���<�Z8ҧA�����j߃)w7$kV��{�Xk)���5/��\��;���ʦ7~�`�/�:\("%�� E	nn\�E["�zu����~)��`�C�۷�-����?������4Ú�o��s�xth��]��^�-��hi?d�����Z�t�5�mUd�e�[$+��7�,� G�F�g*���pc�6'L�[�=T���F̦W?j���7cԡ��zJ�}�RG~�5��:ܴ������1��戭��+S�T�v��n))K��p|ь��AⰂ ���p�p�8S�*���7mw��6�U6�4�6b,H{SU�wBt7Y��*��P4 �u�k�?�����3��s\5��@t��lCT!a�`�R��c��=-���sѡ��񗭅�g���_�`���1���M>Δ�C#(���?�D6�F_=��ٗ��)���'�5K��|��+��;� Q��4���	&�E�dfmM����x�@��H���|�8�;n��.4.�0���.���&,�-�x���L���N���x>��~c]���*�Q2p���2t�4G��ˎ�q#y�5[����[+"��4��I
So���9�4�%������**�(�z �R�Wwg|���v7��}-�j�Z*�_|�7���#�ج0W�����U�~k����\H�Z�@NIL#�ZWH��%�����b���H���c2(bGAv��#����$D�D��n���z��Ǳ�%t�N�N�'��zc��K-$/��	0�m���Zhቋf1��� v��ؐ�}$��p�_���>!�QR���FM�a1�3���RMa��Y0q�)G\��y�8U����"C�FX�W-��/F�B��-/4��R�Ũ����2Ў�[�K�q.�����->�d�I���9*��.��cPk�T]��m��c��B��K '��E�"X#��"������j$� ;�1��Ǹ���'E��ƛ��$z��k�V0�=�l�[ 6죐Q�\n���TV�[O��y�W6qp2x�b��9-)�]�XG�7��_7'�[������5*��Ζ�sa��ڎ!����;�mG<�!]6���|�@���~� �6�$/j ��-Ɍ�����Tz�3�6A�T���L�>-^�F�Z@�mbB�=9����������0�,��y�W9Z�U.w���>)���E�$hoZ��k��A!�!�[���E�a��\�ҫ���~V���<���?8�� V���T�w]����c�e��/����W�M��:&��L:)�6!Ō@�{��?O匇g���KW�-���P� � n]��y�ݏ�e��*1������<	�w�6������T�= 
�:����S��ԗS�U�q�ej:�f�[]Gr����R� 2~��~w��Ɨ�x�X�t�SD��_av��uv#��n��0�/R�=�uE�=���<���T!�J>��������S��6�"/-GꜾ���=�:�dz���l�v�T�!�XN��e�A?������Y�H����ܾ^�Sq�M��ďVj(��A;]K��c�D=m���(m�e�cQ'�^bJ�V��-nl����������w)T-T㩑�!�dN������/��	F���	�!YV��<!�wy0[t�0{�L%��A͝
%T�Tź:����cP����>�.F
T�a�.����������f��mDnL�c�2���*#`�q��pF����B1�ZJD�kY��	R2(���̓~� ����*�����c� +�*�f��*B��8?`4(��kOjk)�C;���{ǒ�HGjw�G��˞��? M��]^oBEypl;iv����>�v;��{�sc�fɷ�������Z�n����^�����S�m$N4%tC�P][ض�xX&\�T�����p���-?�E�����F�}uS�'_����p��?e���Cu�<N�R��<����~`oC�£^%^���M�ؘ4Ư�]QQ�K�XJ��Q�����Vk��n�q�KQ��y��?	�����n|,�
�1�X�����l¨�]s�� S����ߵ�ZX�e=��$�;�e��;uqV����&����|�R�=@��`v,����O�ޅ�1��4���QL�t�����M�{������:���_$�~xw��)u/1Ǐ���o�G��"ӳ���K��5��*'������;*J�,�#[�
8�<;�z� ��|�\��\Xy�Ϯ�D���<��$�kXPN�/��|�|Y�\Sd�j�7�nz_)���h���x"�nH��Ot�d��dO'�{2�c��:=�X�<6�-xǁ>��V�����G��n��Uc�-�"�y|4�:'1��u]M�J�{vgwn���YZ��d���kPB�C���O�N������������\7;
s�Eu㚅�@��~�P[�^����x����+Ԝ,��8A�P�MC7������7�;�d��V��,"�]��������%�d��	+2��\�?v ���!��2\��F�Պ����T��m4��4�/(^Z�7�R���S	��� ,������:1��ݵkM����� rv�	�K�$:@ .#̔!v	��M��2�J���X�sR웪@���N��DƳ�燦��G��8b����u���SPg���.zŤ��i|�us��y�&�yj��a>!�C�[�-P�x�<c&�H���o59̽ݤF��!U����`�tF�i��9:�<�N�*���~Lf�����a������|�3�*>�[�i���=F�5��i�/̏(���������l?�̪��6���r��ϔ����2b�xeh c��°� �ʑ봺Y�{��5�� ���x��m����R�!�땪��6��⧾�H���/@
&��X������e} �4zm� !�����My��{��wFb=���%�u!�X���L';��`��-��a�5��}�� �s�&�4C��N��F⬕��eN�-	�G�㔏Kj2���t����?�y�y	UvP�p7��*Ox|��ce�W�B�G�Z����A��%g���lO&�x⽧��0��m{�=��B���UL�6߀H�ZfR��:O6ά�%͸���������o,D���������Zo{@�l��\nAQ����e����V:V��-� ���ؤ��,�XKaZ[���M�5LE�|�:f�Y���`�9�Hq?�Q%�f�nK�pyJ(2�A/��f��b��ߧ7&H�:����w�U�sᾧ0�I�ߺ������ӄ���(ҏ[u�BE������d�]Ul�����9���W�Q�F�r����u'4d�M��{MYu44���cĴr�!V�� �L0xd���mP<s���~&�Y����#���	�թՙ)DRC<��"�\"��Hד�cV��5��V��U}��;�e]��{!��]�ֲ�VZ��T 9H�Uv���7���c~�k�3Z�
�+f?h�\�z����N�ë��s_�.� h!�ض8"�|>L����m�է�Uµ4�E�AŎ�90K(�ԟAiTPO}��x6���VpHԎ��&Ϊ�Q�	�����QV��Q�|��P�!ݤ������9��
��Ta��Nh�w����d��ˊ��N��)�V��F{����F��`�81��q�]iP���f��,����q�I��l2׃�݇���:��='��;�j����	��f���6�r�PP@A~>���3
�)E�q$Z��E�<��DF�R�������r��P�-m4���;.^T��|�,S�࢖�Иj�q�_0���Q�\�#(Hk;c�9��l��.�Ѩr� ���:�k���.ʶ��;��Bv��S�|�c㾄,+u!sk�l�@+���{�&��0S��p��a�?��h�I�8F�U+UN˵ Mx=!���+����4��;͌��P��b|�|\��/�'�!B�fD�����U�{�k�sW�(��t�����xWͷ"��Hʅ���;�O�w��h�~;C����Uw�3 ���)�7%��2�z4k��;=6Z��V��h
�+B5�T�H��ڲ����)̞��@Ԓ��B��D"�z�%%YE�L��1�*�U��d��ar�� V��;��K����؎W��;?H
>bC�i|���۴ ���)Ԑ@/���������O�$��P4]�*f�*�P)�?���v���)���]�� &��$C���
����{t�	%�I�<� ?gC�&�<+��2�{)��Q�X;HNv�Wa��� F�*td�d?�7]b���?}=�`(��84p��b)�;i|�A�'U5;�HM��/�s��~".�3�v��"oKn!O+�uus��5�R�������kț�@Hp/��p@�W�A�l��d��Ol�k���?���f����wˆ:�hl�]�l3=5Pgbٳ��%�;���#�`Ւ���y����oGW��q�ܺ�y���^�����/q�a������t-�,}���@x��P�(�_3*I쮌�F�����#"���0���9��wj���_C�����o�4�L�D.�ZT��?��h�G��j��T�$��(�X?���ƴ��n2����']{��u�8����V���C(�OD3{�us-]��� ��jB�9=b��a}8S��;�;�m�m3V�ĭ������ţ�Lj��]H��{�K/�!/҄���Ko#���=�P�[cO�k�j��_�E~�p��6۾�����ȈEG�ֹ-�	FYa���t��6^�t �/�o�����#�-gkY�t,��h��Ε�A����7ԪK]��т&=}+�4���4%�1z��N�-`}ѿ�{^[�ɝ�z���j���=]q�M�Y8S/mnz�a��⬌Y�d�S���_�-��M�̱?6a�ss�%�|I;�k{��.�r�,�x��f�W�s'���=�j�?ЊJ�3�HMK�%dQd�F��!�ȍ)##p��wۃ�:���y6+�OY�_!��q�aLAáv��e�.����.+[d[�A�A�h�J��N3��!��&���1A����Fǧ�(��Q����f�/s�.�Xx�"z�O�Ԙf��k��N:�׫N�{�	(��5��c�~�W4Yԉ�����ԝ�����!�'i��'�;j]AI�H�����g�&��k�_�e����8V'"����;w$O�ͳ�~3`<�˿���宎J��â��gF1)Bė�ϖW|�������?���4����a��iԨ����z�yN|��4��>����/x�+��u��������9u�,�/̚�Ux����9� g��c�A��煢)���3ܩW�j�p���{jV6���!-T�0�`z㶅<�
���(�!TB��iBY~xEJEA�V��-c��n
Cl"B���Cad���k��넾u�_���i>�K3�X�jZ�~^f��M��:�K��`W��ٕ��uLzM5�W�1��� �BJ������_�"O�N�T�ښ��!��R݇܎��F�(q�p��\�E��P����N����>�j�Zlf
Ň#TjlI_�[f�5!�e;�o���,����$�S�%��g$����j�|�$��9�f���6"D'���w)Y�'�!>f�����'���	����"�aጝ1"fW��X���e�f7l0���=��ti���$\ ���g�¡�w���b9�#�Zp�����Sc���x	�O��C��g{;�����AX��7IhK�u����-��1����x�_Y�E�+n�E�Lj���O�����jt(�e�},f�l(�)����=��;���hoԔ��=Z"�g=X׸i�xڛ���]�~���J?�1;�q�j�/�dE�!���x�K�Fe3�#�}S���F�;��(s,��I��Р.��$�9S5�|M/��{^=�Dg¹P<ܻ,�ƌ��F����R�Ε��t��e�Aך  4ٴ���X ���|�T�
A���	
��u=���8x�O��0н�R�o�X7{�-��]�."�C{�Q���E[�H��0��A@U�ʿ�7`=&i��=��ִv��|���=��g� �[��F��t�Y�)0��1�}g�z3e��K省wkB�jq<Z�h �\���\s)[��mZԋ5�ڇܡ�:`� ��|�1�����_$��2��*B~����d�~�WC��뗷lҰ��u��!�H{r���v��<?9��-��|Y)�vX�U��Y��t��An J]^ɖ>%~�j�).�oP5�.u�����s����+5������N������Խ�dܕb�(�c�a�`�ȿ� �=�K�$ж�#�Ly��Zy��' tv����f�Ao/r�b�
)��e���$�d�r�VA�Hu��fa+��|,&d�ׁ�3YOdf�|����5�%����H+֒s֜v���Xj�"W�����J�Nׯ��(�,)�Ȭ���m�C��V��6_���5ZC���`n����9�1tk��^Kj+1|���{F�n�Ҽ��j(�/~Ě�M�����cpљ#�
�?��P�r
ህ�em�D<0�5F��<C+@�{f쁹.G��k�������)L���b�î�Ho��y�e�i��G���a��5Hb��!�=���q�dq�$׵��
��򪭯,ԯ�Mzf��aN�ޔJ	�t!�fyS���*���f(H��
۬��h.a�)䪹[��I��_|��V��~i2�:0a���(�NΪ�B	{Εd��v�2��zGS(Rt��g^�o3}D���Aq�H���}��t�RP�����0�«��Huڈ;���*�Ȟ�O\K��W0�=~˝��P�wſY�p�/������=��մN���y��!~�<'�1�XY�+�ɨp�x��ń�����8ܓ�:��8��9��d%�.s��~�q��n�fϓ���5f9!Խ�}q�;g��0z�C�}n���q��&��Nh�%:$X����%4�A��7^?j��P�d#/�B�~�,t���̺����f.8���џ[$���<W@��z (Z<�ko?��qt�n��=gW9U���VT�p��.q�M"��D
�n�TE
t}Z�Y�>�f��>X���8/�9<\�^E��ד)ƪ�}Lɉm�RMt�,m������e̉:�l�v4Vg=�r�s�.ϔ���f�z��)�cբ@2���ya�ނ���}���)^�Na���\��Z '��(���F���.�kx$�W0*��������}�KuDG��%}�-��ӚNi6�u`�}F�A֟~����f�-q��Ůs����-(�)����s�.�Ɏ$��[�x��rk��#b���mϲ�WY^��Sy�,�ZɎ�|�a��ƙ6�B�cJa[;�v�̅�r����|5�#�71I���G�A�8B����b�3#���������l��: 3�0\��"X6!�p����5�[�P[�4#��"���tM�h&"���u��t�y�,�P�����ڏ%qG@��Q���c�Źa-i�ƒ�Y�^��Ȩ��@:Xi�"�:7��M^����?���{�y,vEKkl�����ƒ����mB;͆�q��-����54X�-@A�д�l�^��u�'�<"��B� ��n����A�3\
!��)�����)��H
�u�4���Q�|�ԈI�ٙ�!jEL��/G�=�w�{5�D�/U�=w�dĮ{��IH���9SM-vϵfcn���CH��_
^��6Ѩ��U.!6��.j�H2{ɮ�2���QA���0?)�2�J�Mg~	n��w����i������%B+���g�}\�
F_n�([�tr��g�m��*-�:1�}fwy`�Ϥ�oYQ�D(��hE�`݄��F�ic���.).��ƨ?�ε�R�>�^��Q��e�pJL�!L`�@��>+��7�o��<P��}f@$t�]�5�/z�J�����yZ�LG�A_�Bn;��-�rVW^�m�,���)lmF��������Az|p�/8��Hm��J�s�Y�x^��=wR��V���^F�u�5������l�pF�͑~)��� 0���T��#2Y�[��ݕGKK�9�_�0vi�[R�@�V�_D?���P	��tM/��b/��&#ތ۫K�"����(xAH�C�4�@׌f?�N[n&�M<��8�[�}�-E��$C8�d�F��kBe�[[��W����Ɓ�@~��}	�'�s�j"'\Q/wM�3��<���C
�ا��G�i���wq7v���vB�U�O���D9]R�=���3�r�uj�ŕI�.#�W�o�h8��?�^�v�{Ml±���/�P�2�%$��av�T�J{p���OG(A�W�6
�Q �[�G<�"	�β�W����$I]�m�q~���j����������w�)�_(���0k5c��<α5���)�Q�Up0�qѹ��;#g:H�2ˤk�@��Y��==������::��v�ԛ�^��{����	�� �P�yL�L])8��b.9�w/�����*�K�	��#o纲ضL%X���᪦(m7)4,'/�&�-�j���ݣ��1��ې�+B�r(�1�<r;���xr(P6N렵���qRa�U��f�U|k<�As����A�[��;��n��&�Y�'�Ĭ�}��Y�$ Fy;m�c���aTD�NxO��;B&��Q�ƫ^���yȀ��y��Iڢ�^�'>acW}���Z��A��$T���$��3W����0��<��d7�u_p~)���d�T�E�.T�܏[(�WdBg^-�'�i�iF2�߶=w]s�+�3��o����61�.�*<.2���iQ?Ԓ��6��]�tU��3u���}Qu��+�l2S+�!Q��8�,)Le9�exH@���*?�FZw�K�����U&�Z��bi��vnq�V��Q�b^9����*����_�_�e]�9��SU-pژ�;w��*�OM�,K�pG���p�'$���薫�<d0�ͰQK��`�)��-n�FƮ�鐌۔)���6?�c����;��1�6
z��w��C���f�-���a�<�T�Գ{�!{Y�Xs��I�.�U��(��@�WocMap����"47�B��'��Q�:�P��4�T�z@�����2�h�Hk'B��r櫷�@K�K��z�lX\�>N�hkЬTwǅHh�1g�a%�À3PA� i�v����P�b�Ӊ���DQ5l��2�+sr�b�r�
y���L���w�x���ܖ�c-�o�h��z��<�O���٢������֤XD����O}���UU�E�2u^�:��{�/�f�J�P�ꖔ����EF8�&Q\�|�Yo�˳+u�1|��=D[�CWpx�j4���B@#�C�G�s��j�����8�$	:�2��G��7�T�H�U$>)�%���"Zg�FM������jG�F@��JX����}���"�x�'��8����GO�ș��XFNɋ��U�o�0}ْ�j�q�h��k�]�ϼ�4�[��B�q��Xw�)�1$����2U}; e�N_�qr�9b��˭5��a��]�WuJ��ٷ5�䥠���Aʏ������MC����3�уk�ܝ��q���g���ȝ��f>�[@�D!�b�G��$�ocME^�T��ߪ�+x�����������^��zX�<�/0��4I<SK��O�eơ����l5�
�v�����C`�2)f%-����3�������QGu��z9��:?T}ʷpl������倾�!;�i���10]��Ƌ�&3k=���Q���N+��Kz�+yx+�GF� �Tisg�s�@T,A��&�����&�iא�,tJW^��<x̊Y*6U��͈����(s/�e�b�I�s��O�ҁ��F�;Sߝ�鿳b�U d賣�b0��<�1�����H}�$s,:�F�
���ȕr8�I�wl��c|J{��d�b��-��|���9�r�� ����bfW��F�o�ye��.;A�B�������1!��Q(�FK$~�kV.�Xӎ�B?F��d�t�Oh�� f���@V4!w@b[����9\�)q�ay���5�,��T���8������Sh��r�ӵ���������>6��g��3�l���g�ALq�Q�X�fH���5�JM���-uem��s4�{�I��@��.̫|��z��8`=[��h �Տ*ӆ��U�P�Ҙ�,���Y��s���4�c��Ţ�l��n�?�;8_��bq��:$(�g,	`	�o��+o4,+g9�����uw�`�t��k�,��&HK�=���"�T_k�.�$����V�\Ҝoq�V�Sr�OK���x RR�6�	��f����Vu"�"�*��b� ��1�P0D������'M���Kh`�vc�Ө��Ń��q!�2�N$��N�%���0!�+hE�8|��-���$#ڄ����·S��R}a����(�^���[��<6҅-�!�?P�ў���Ҩ��^G���L�9yKm#OK�Ff��BT8�}�b�D���Q������ .�U�9� �x�Z�.�3��Ϣҳ��\1!��%\m���vC�@)Z�i� b-<W;'
$3#[=U���VM�#�>|r�7���~;z�6͊.����K��N\����3TxQ):w��%�Kd��A������M������H�H~������09%I�w<�ւ饴�AA������"0츲צd�h������ ��S?F�3�������y�����НC@Ӝ2���i�@	��y�E��H#i:�ٗ���Tq��TV�yp���5�M�E���3��=�tf��&*�A���RdCH�q�A|�]E߱�����({f�Z���!j=����O���*�HT�Li�; \����H+��b�3�
aS3`�F噎F���/x�h�;z��'�ىǟ�H��w�B+�>NجDS(�}/"�5��&d��T�ǋ:��{L[-穄����gpϗ��D��K����_ȷ� �b���1iM�N�P?GҘZ��j�o+ԍ+?gBV��BuZ*�_{k*��I��)����6���TK�$x�|jL*���ǀ��.i-sZ��=5*�X4c����|�t$(bs�y`B�&�|ZB���h��X��f�X��D&���]g�r퓑�v�����|*\�_�J0&��Z��d��C��f�3��=w�Tz�a)����)\�R�<��l4���3��0��;=���V*�u�'���b�	�ݤ~���x(���F~��#�,&6�����N���3�F l�졕ٖ,;�<����r�)��g�q��W�p[
���v`��20�Z5���s�J##GiM�ps���l�J$��D�~���W�0��]%c�4���%�ׇ�	�����8h��y՟����P�:�%@�E}f��=9��4��PF*��(��V��6�p�CEt����.
�$�?
�^��ʹ�|P0�TbK�O�v��GUQ&��s�3�W|��Nc�wt%'x�Z:����zs�'_�8�3��&W�E���T���]B7ؓ��2U�Kp<����G���a�r��l]�0�4,E����Y�X_�q,8o�8Qd�������X?�����'7�~�(���_�_�<��L͡�?�.����a
��b�ٳ�r�-��T�ݼh���o/��@?�fE���G��p,c�H�uxж���z�����-���iu�ch��
�ΉD~W@@t�8l���'ր�;��7I���u_�{���c�	��hr�L�-μ��|ԖLH���*Ya�v`�E��0xj�!��6NK8����x{���]|�gOHde���<��ާ��u�n7!��i$��q��"��N�E����/�]*�l���	dv
m�o"�j��I�Z��>t�����K��d�l�r���(zw�����i����Y×%���1���%L=%�O��Y(g]�EOD�M\5��}i}�6����(��H���D�۳r�-)�-��1ԟ~�8�]���3P��}�l�m[y�!��0�_��	C>��P�@c�\s�o6q��5���աp��R:O��v�\��;�4�@M+����H�c�0q�Ỵ�Y!ǚ�p���;�+K�+���fr81��N߇���9Mb��i��Wo�)<"�_�$��I������ @���.I\P����w�kո�h� qM(F\9�<^�jÆ ���f�sNy���A9lմBv�mZ��ca�T���PM�v"0�NҌK��7�R"wU?��/3����`�Ѥ�eK|��I~��j�)~�Z�j���.�M�e}&����f
��+��0�ig�n5��@�������9���ν�.�@K���q�>�\?���_�
/���k�uŇ4/�Lb���Ʃ$��.���������i}7.h"�����J��.C�6+�7nU&���
�z�f\ƈ�R�E���j�<� +�aG��Ņ�S����&oM���qo�K����@.�p��*�`�4�dCh���~9����)�/j�0EE	�ӗ�iELY'jR|��_p6|��\P�I1��r�-3�k��*��?KC�D��ny�N�FL��@ �X�5��=AV���WaN��N��h��C	��z�oS����<J	�M�$cR:��l�'��D��/B���/�*7{r�h* I�gIt<��j�ۋ��5�?��
iR�.7߸�.�AD@Cw��t��]�M0�G����WEJ�a�)=3Trv�]�a�Q�4ہ�3R=q�`�i_��n j���ܽ�����LN�0F�����f~o�^�h�;4ƽuMv����j9y�*����S�&!i��T" f���
��\�p{N�$�:kQ�������J�e5��r��0ϚRۋ�T���Vh{��[฻3T��4#�����*� 8���'�Y�~�>+�d&*6nL�>Y�ցd��Ȥ��Gy1���&�����-��Ud@�(R$q���oc�9�� ��4ta�p3�RI���Əȑ2/:���.#�*K`]��Tд\ �v�
��6�iۃ���ȣZ���T>�
i@���;R�ψ�.]Z�
[��5L
�;�򥃛9��	E����9GsP �iK������R��v�`Pξf�v}��େzsȷhO�� �X�SvC?zr�2*�!FhB/���`���<�8#���K8"l C���U:M�ہ]
�O�G.9dPc�ݐ�/��MP�-IA0�bN���=��+�P+�o�VD���&�*��4����3�lD�i@���c��#j$�%�
N�aaˣ�>�qkMI�<�g�=�܎�'ط$�V�e]���߇3��-
��Q:�.�*l��u�c�_�(�i���rK�)gbmb��=کy��b^a��z^Q��t �����_h��ө�q�y�SB�������dQ��=�|a�В��Ʈ�����}�3��Q��Yr���x)a+�����b{�g��P/�.��*l���_��J�rM��|��d���g�og{�D�<1��m�<�	��	��l�����{�b�*��TUM�Tޔ3yJr�aߣ���~�ښ�[v�{�@^^R.����� sAh,-^1��#��GP�D�1� ��jsalN�Q�eE՝.��Z@L2:?�9�)��;����FD_�hv3�4�.���+�@�>~[U����O=�;�jR�`�)�y��P�1��+�n@a�{�T��q���p������>�����N`��u��}&�����A�(� ��8QZ~e��ِS�b����\���5��]a�:�CJ\�^Z�"
¸4���=PZe}!6����t�d��a@��rda�W��L[Ʋ�(����_��;{ڽe#�tV��������/��ج��t�
ŝn�{�XYMC�vB�{���?�R��r �������e �V8eAO���Tuc�U_ڈ��!��1�=�����>�>=������W�SV+ْ?���P��%�m �&Ax�|�l����9\o�����-ſ�2��\Gg�j]?�4	���t�fΧN���A�~�_Ԃ���˂�j��}�m#��6\���U �"�.�#0!��i��6����"����,�VQ�<9#�3	PX���j6���0�lh���Iq(r���2��w�z)�g	�TA�0.Q��հ���f8bF�:��.���typ���a���rV�n������f+j^�ʡ����z�kw�+� 	��EiIKO�O��=�����
��0��J�.���Vi��>�z#�:�^ �'Ӈz/(2�����"`:�)��7�rJ��xȦ�����ͼ�'�!{�H��5�L|�D�#���FwF��f=:��ұ����r�߀��,���E�uxݫp�G��2_TLv２RuY%>���'�,�#/�-)�Ȧgd�# B%18�Ï0�������l[u�}7Q��ߪ��u���(;�N�v�a1���D}���w�<��{QL�{�U�샰���28a'd5�~��"��f}:���I|H8-�>X+���Q�r�V�g	�Yt�kѣ�Sĩ�, �%�vwǩ��f9��i�)�}�찥`�'���Z~5r�}u�=�]Sl���YU��Clɔ����F>(�Y��u�a���h��P����c����4��eIv'&�;��9�=�Q��G�7��.�r��ݷ��1x;��t[�p�l~���X�����P�u�dq�9O����S��V�w��j��kr@S�!�a�"Ѻ����v����_�1�~�иqez��ٌ�|%/����P9��v�����F���<��O���4�$j��$���:H�)_���h������;Z���*�1SuE#{��ԸO�v���`�f+�����
��b���G��������&D�:ӠAGh��]ǞV�8������>�eG�^(�P��qQIX̨���F�x-�H�<�A�:��nQ��
^�\��S�{� ����&�b�ehTR�g�D^;��,b�n��7u��ɑ����3˘����f�O���گ;Jۜ|z�;�Ԕ����^h�I�vE;׻`9XV��0D?�_!����wٖ�7s����	�+pBgm�Y����!Q\-lm �J
�oU��������i9�C�W�" o~��i�`�����l�|z�< 枳�C�n�r��_[^3�c'����mj(�'ئ�:�|�y_
I�ɀ��|n�w�=@ї�Zo߻�sW`oi��D-��Dzkӽl���I������S(SȆ&[8	Ũߜ,]�i��F�n.~=�Z��8��"XBH"�˭ (hr�P��o��yZE����b��͡���ʻ4J�ǧ�H,�0�o��윉��V'�~~Թ^Hn�O�}���dԙR��0��L��f1W���B�
�%�t�;�V������USv�@��oE�����UXw~�6 
���1Ά9T�v�nGb��N�K�T�(|ռ�E�z:��X�U@ZDԩ�I�gV)��N�WieS�a� hV����EyB���i9�ko'(xX��=�� ��?>+���V��9�]x��ai!]���bRwhQ��0�6o�4�t�9B�r7���j�7����a�}E2�WB�Q��!g�媉Ѣ�kkc��洯N֬�3Y\>-�Ι��41�mo�RP���s�
&8��?*��ƌ=�5�7t�G^������ݘ;�"�E��s�Vj_ܽ�x��d[��?F�F�+/��ڹ*s���J��~]��{+�혘� ��~
�R)�4�	A�[�	j]�'a����x�A�Y�:"'�u�,�Cm�E0T��c_]@�B�*ـ��`������?%�|������e.Iq~�N���	��x�@�����U�'���<%���';m�mD�B'(.z�('�IV�3��������O,4�g���5(�j�L�&���l$�]p@`%��W�݆Q�2��ȋ{<�?Rd�D}$�>='����br=�L˲s�I�mڠ���QđPvs&��+�$٠[�'
�=�s�b�{���`�o��D�Hg�m�S��S��!e�.y�R�nXl���g��y-J��3db��e�I��r�� ��hJ���|�-�8bg*O"��(�֡������!}��	��1����N�gQXk�ː�-K	�Fm9ׂn�>�r��_<!��4��bĜ(��J���*q]'�?L�G��S�qfq����"'L�Ԝ���X!�����m#e��9�LcmJ)\��Y�����+�mm�4w��ZQ\<�K��U����i���iu� �Yb���Ǡ�����n%P�O�9��h!<��}ļ���;��K|"Iu�+�M�q1�Y����>�'��	?Q�:�>C��;>�z��&�"�s�@�߆J�C�����tSC����.p����c�TƔ}H�MݼL�����\r���kW?`�D�d�nm���*�ڿf̚����@<CM$g�Z�gG��`����t`����]��g�V(g��d�i=��L�*�F���Lw-<C]U�#��l`���i|�T5�4{�J(��A��O]��ǩ�/���|�Nb �j�	pE'tڝ��*b��?���'�޳y�92�Q����j��X~�|_?$�ݺ�d�	(l6�4�^��I��\�zqJ�3$�Gձ	���Չ��b�â�K3��TRh8�����4,�F<�RK��в�����Z�׀��v����������ط�H�TvpX�h�VMZ�{T�v����,���Uc$�^��qm2��M,U�+Jۑ.rAw!�9��2��9����n�"��I>�[�߂t��`�c�-�̠L�+�6;�ą��E��v��IA�w��o�7����{��̸��r�>Z[���i���S�;������(5
��򀅼z�`�k�F`Q ��K����Z�J�ׁ���BD�G�\��ua�>p�Q�U3j�%R4ު��vF��1~�� &H60΢eY�<�֧�2c���;��
$d�qԔ��QMNe/n 1�V�������7�����ѯ�/I�_iƃ�L�v^�:�O�O�*G�*p������� �mUb/v���p��	�=b�<K\�5�7i>���@���%JHL/��b��������()i@he3���������*G�nB��uf�A�g�'v̳��Bsz���Z��2��V�,3�!b�h��iE���\l(��w ���v5V�_���oM���J��#]nAc͞���\�9�sЍ�z���j�#�� p繸�b��e�v!���8�{f~�_^��e�l�r�)�J���
�ƪ�e߆\�{��!�v�D+�*y0��*K��$�=�z#.�%.��5j_������F3l�U���_j���P�5=�|�9�=�4��m���;2��r,n;h����AI�I�so�-��K���b��'��T!��RK� ��#NȻ0�,����#�j��UИ�P����V�݀�A6~��w2��E��MX�9nj��5!�mp����i�C�*2��� ��D�����`�M�Ø������@O��NO2ҡ<ؑ��rj�����G e"7��1d&�6)qkh�]?���I� j��Q���]wr����|X%�d��A�~W��u)v�n8�D��˔�DH�_yk)4����Fޚ���Տ`�a"Xeb�r��[^n���u�4�V,��a��L�g�2EJ�깺>��(�t�kܜ<���R]%�>�'#���C��1�|_�G��Qa��[%lO���,>n�v�[�3҂N��-o+w_��� ]�w^�<Ʒy+�c�V����r�.���2���	�PleLgn���k����A�j�d7���9Ol��!�u�dfz⻈L%޾?M|���t��"�'!?��x�?��
{u�ygs����^��-V��D{e������a��F򊙆X��q��S΍�7�a,�qDY���ڄN�7Y�-��܄R0Q���`|���f����n��e�򪯎P���(?�cLZ�{o��Ԥ��(dFS���ߙ��Ii]`-a����5=*B�_��vp��JN���>�)�|��Q~���^�2Odc/p��� ]�Y�� <r��������W��~Ҩ�XB ������)��D3�)����.�a�f�	8V�݁Wn�A[.t�|�l�6E���w��@�\���
F6���h�JF����z�!��k�Z�n��]�>5�nf�>�e�xМ�YgU�k�r�K��\�q��6��Sc=E�!�}Gߍq̓P (��o�vh:�"�o ���*����SKBG�q�F��c��4�4��;�O����R9�G|D��+�R7��0H�݃0��j��s��{kd
�al��g�"�mz�	�R6����*kh;�1�ozC��鄊B!��|�H��P-�3Nt>��Ri���}��7U&�q���?�H�� ����Κk>��v�cj�΄�0�/LV�䝎~�[?��	�A�&��x�{H��<e��lM�5�/�>GBt��2�� t�2���������zGOߋ�L�չ���V6k�z�`�Z\�͛�yg�(�%��� RЇ=�A�`�5KNŸ�|9��i���H��#�,&�C+�����k���HM��C�*��R���Gw2�j( ރ�dC#c܌](X?�(q�TQ��˴�o˳}�Ns���~�*�)�/�I���Ty��NV9�c���2,�E�if��=d��f�}ܗk%����|��
�v$���2�ĩ���n��E	�G9���K�����w`��1�l�֢��?ɣ�~�ZBc�i�ppuz:���nhyS�>A��L��˒��!{\9+���2���Et_�ǣyJ��޿WQl����l�y�E��B�=��N0�us$o��V1B%����F5]�cj��q2�af��Z��~ك䈂������fv���ҟ�X��R�.,0��./����N����O�c�W���BR��s��0y d�v�8B������ἍdmjyK�w]lԲ���ͩ�<y���;�6�ך��Y�M����
\�v�a�3~��F��'�|�u�%�Pw�j�'�p��2M��o[c�xɺ�'C,�O����<��j��;h�SA�p�i��:�Hv����hC�%�&ƊS5��#"q�6J�,"���顾<�Jk0d�����o抅�#U+\�n�kmCT���y0���RA�d�ߘ5�����U�����،̩ޖ�e�y�X!K	�Uփ���U�㗺9�[��ץ��������q�����w�|z"������@ϒ(=26��!{*�ܶ0�3���kq�95�yz�����&���U?��E�U��$�e���.
�U��}{��u�G��UCy޿�4�\ �^!����]t}����������Ot]��������I�8nO:�f; �m��Pd����P���d:`�K1-��U�E�Vp��r�)U����5x����Sk8��Zb��;Z)(c�
�'84b��v旑���O��syּ{E�Y��Fn9W�9��Jߺ<i�sX0���	SNR��Z��'C`���1тM14VW�4��Rp������(�&��ܓ7>�02�u�O��@+ZA<�9��� %�Mx��c6m�_���z�u�hk6�L;�nj��C���+@;�Ц6���ϾA
���8�I�C�����W˛Xe�5��J�fR�.=�Hݦ+��+�S;�N�+���vJ�d��p��O��Wz�7wȄ���~�	�V��l���a%����uN}>�x'uI)<���9���1P�"lE�bbv��L।�ԩ(�\x�v({���ܽ�b p̕�",r�j�5�R�@�������>����;�����zOiƌ����a��+ʗ�;����˛+��
���N�V���g�?��5A�44G����is��zZ�ɷ�0�?��L^��+-�b�۵��
�HaG��M Nx��_A���,P
UBP�]E���7�o���_=F��^m�ٮ��sB ����OD%@k5]���� \���WW�q����?�5S$�����W�<o�������q��p�\q�m2�9�(�����������sU�]F=H^�/m���C����_1𮣴��0b��tQa�K-%@w�����V@!,�~���
t��8��I0��-(�E%U!�q�e��/�:V��3^6y'�g����Md��w�)o$�=9�+��i��U-�M�kk��h7~�`~Y��E�״78<��46œ���u G�|�ћ�V��>n�&|m��QX�P��?O���H�e��M���]�hkt�Dg��=1�..TQY�����O����n�B�/��?�Wl�zV��{��Wb�Qq\Ơ^BÍk%E0�a�-�/{�&�
�.�a0���� 7�$y=�X:d�"��;)]��8��؉����(#���u&c�h�4�a��n�1�|�ӳ����E6l�)�9�Vk�d�E�+����ؤ ����`��Zy � x������M���+#��m�D��}��~�ʠ���v�Mn�p)��^3� }~]^�5J��{�13 C�/F��-�1O�hZ�6,��Ȝ ���V��p����15�$�>K��C�N���zO�(����}�A�Zϻf��g��*�g��,�R/�E�Nc
oL�^܅εV����y���0á;�05�W�FO���-���Ǘ�:�Mk{E�DU���� +��hN��o�18:�A����[�R���Mˬ��&�!Zv�b�ֽ�^~ 2�;�Z�ۏl��1H�,n�О�AĹb�'��Z��a�-C�o�5&K�:-���3@�L;�l9QgJCbA��g���<�Y��V'��{L��U������:�٣Ɲ�V%7�]˫jak>k����շ�C�yOIrnW[�=eh?)�AV)O�(��BL� E3��<���݇p#P��Fq��Y=`LT���F�q�%ݱ&P��WY��c����(�<"Q��<{So}�6m.Ih�#�(��p��%��d����4�� 5��.�݁M�����JW�D���A��X�`����p;���\�ߗ�a�]���~I�5(a���>0#%�
��rX�6�1A-q*�s�.�;���8!���	�U;����� wY�@l�eMlaJ�����oq�2c���?縡N��W�1��1�����\S�m2џ3�Ļ�侃��j���#��Z���Ї��k�E�3��3��bA�\�7���t���	F��}�48���YT���8�Y	�����nD禅��AE���hw��at�`Pݩ�ɭqpy_8@&�3u��Ę��E����P��o��3���5�a��pC�V/��S6Sۗ���<pW �7F�iD_�Q *�+�������z`�n�k�Q��d�h;k �zk�MJT�f�PA�Ǐ�n���!I�|;0� z|Ɖq��f����c�"'Q��˭3��U��(���kN����Ւ�dzOn&T�e�{����l��J)�8$�������k�:�r��:�e�.Θ����/<B*n
�am>
P; �F��2�Ns�3��E�I3Қl����u�h�4+�>�_0�6���#��� �ai��N��r�w}{8)H��5��w�g�x�6����V�q�CƟo-���;ᱷ�� � � �d}wXw�X/SpCZ�je�#�JV3H���Ww�Z�T�� cYw*͢��s�����R� +R����ĸC���a����}��b����u�
��ң^_o��?t�&͌F�B~����@�N;��U*�L�9���[�w�w�L��>'g���u(������B/���W��1���n��b�����u<׊�ʺ_�H����D1-�?�3vͮ>K���'yhN��:�!�l��]�Ԛ�����G����E�3�	-���M0fDE?x6M'�H}̠�ƺQ�Q�V�5;f���+ I�	��

�s5�łЀQ~��T_T�|�̠ɍ����YEn�']��ީ�=�>_�L�6ÿ�~�BR�<�����2�l+/Yqn@�{^h+J�!��)M�ۜ�U����z�m���ڐ�b�̕x��9�'_��HC�}wU @�J�Nc��_��b��D�`�!)����=�n^���8G�?�.��J��2f��d�s&�8�P2�Y���ǟ�c�&��SS�;��fA��W�[?\AD�b4|����oI2�p�K��E���i��x[!��ޓ��^�k���N��p������ҁ�_X�n���T��P��QrM�?N^D��/E GX�j|8�݇��Á ���j�y�]�(R҂�D�v�yAY��t1��[ڨ���<����}��U����<��Y���v�'�ʮ]��9`��� ��q����>�H��=�G�:�)k��Qz	��"���$ڰ@i�\Z�r��r<��V�]?��G�Q,�K�p����_'"�R�o
G0x�v��-��si��[5��щ�چ�ؽ�L�*��D9.���.B�i��)�/\ʄe�ϥ�?1)����Tg�R:�T3��/lp�\�{��N��;���W^�a#8&�w�YQ��x�]�s.h�T�V83	���)��o�sh[5� ����|ˆ��,^X%���@�f�$׸��?��<�J)���PIC��1���f�M�"���Q�����.�,�� �=l��`���j��߆ר����`0ܘ39o=���8!C��7������A20jށD��M���|Q�U����A9��	�/��2wb�
j���H��<c^z�!�׊X���P��R��w�QA�,��rO2�������P<(�zN��T�M{8)��g͏��}7��~!�X9��������Zs�PO��埥B�M�r�e*{�ׅ��.O�87�f�|5�����6[���Cg2�de�����~*�����$��H�6�jΩL�(g$F4�+q�=�&����z(����<.�<�� �Z%��QSŗDL�৹�gG>dgg����������A[-�Dv��"[�q�z=��+'ؖG���������T5�� ����G�y��R�����Y����+pN��K	p��n�T�?�l�zA��[�=�l4IZޘ�Y���9��I�C�ڳ[��{�������2���W��~Qw������kM,��j��E=̣�j��>L^!ޡn^��.� �k�4���%wt�7��y/ �@n,�>憕V!�Om���,��h� /��>�mO]��8�7������5��ײa�󎪀�g���چ|a�V�7�ep��i�&�O�ROqj�X���U5�R�'uX�7��I�$q�R�үJf�t�t�H��ȝ*!��åa��?׻�5�A@�.c��F��`�W��!��؆�Eu�����m����R,��|(�%(C.O�B���	H����'�ųC�3��\�c/Β%�TW5-�2 /���3�V�QR��A�A2������RNWE���ِPf��L�$Q�7"�`�%M�P���9m�KVi��?�u<���T%lU�(�}��� �Ǭr$RW�c���ќ����Łj([�grы�F0#i���*\C~��,�mr;�}�d:t�W�0��>"T�Rz�ABD;�o>���`�����R�U't��?�-�љ��J�>X~��Ę��n: +��	k��AVc����w�\��OlJ'�N�]��D��_��� VB�c�A����C0�Vv�t���:J���|`j��� �fU V0�'�u�����K59�F<. ˧��Ȗ���C#7�!�}p�
q�@�.���#)+z�6O�U�bB4����!�E���P������q�Əot�TA��D3Z�C���*�Χ��p"\F�?�0AY�bS�=��7�����A:sW������hx�rɥ�[�7�	��f�Y��������q��VV�
�,���)��4/��2��DB�((�I�w,������q8f��uMݨ=��'��}~��uV�x9]��1F͞�o��)��q"�⶷	W�P�h���`]��ΦzN�K4Ahh>���u���;P��,@4�D���PJ}��U�SJ�ޒ�A�����h?��3�����KW	f�Z�ƈv�MO�:�i�!
��rjV8����5U��ޚ�I,l�
6?�ר�������\)�X� R�3���%��HNѥ���;�m2��hM��J5��ױC�X�n���r�+�w g���}�.������(xJ5��id�3���c��F�?�TIK���C�C�A!̓u��r����G�[$��ּ<��盍ީ�OzI��̬g%��5N��<�`eH]>��7�]2�?3U�7t|I�:�	5���+����HI��BW]:��w�ن|�\�V#�#i���D\)��x���b9O�bm��d��8���l��`�C>��jo�K)�=}@o�Tl֠�>��]i�M�8��Gw:��s��W�ʌ�|�m0\ݖ�R�jZ��w�,��7�)�#Ls�v��r��Q*�h娯�����'�yk�]�{����!i!���X_��I5���v��#����P��m2�1��*UU�*��]J7���
@pp��R�ZCS��X\��Z�Ծ�3��$�Ҟ�Ƿ�4�s3}�Ew���������U�;f�����s:��b䕐�&�����F�퐂i)���hLhj�3��U�"�g����VUF��z����31��k�Ѳ�}�N��R�T2^�uB�E�^��9z�䶇z?�v@M��3�J�C�o ��{�RAU����o͛\�2[�o��8�L�I�����dO���C�už��x�G�>��'��S|�g:���Ǽ�9j�al����Y6`�!��c����c�D�qM���  ���ey�,=��e��1^���x	���ud�]i~�t�_G����y���=�i>z��z�
q���UJ�A��i�<NU�K{�[o�p�����o�y�- [���n4�Ѽ���mwt�B���@��w���SM��a�"��TAx��5�ۖf��)����Ho3�V(��*/^��[�/�k�i#|�#��]�D�i�P�?��FLJ�lC���1o3_ͤ�B��O��Z�5F��W�Ȉ�d��;	_Yo�6_�#�y& �L=�C�7N�w�oF��u�k���F�s"�nU �:'b��e�q
��B�ڃ�<�os��k��c����|Xk��� #P3a]�K�a�Ϗ���#I5Բvq��6�)�Ʀ0�|\�-��h>��������Ȫ�N�8Q�<�H5�J��@��h������D�K�d}��5�������:���2!�
	Yګ:JDR����0S�_�̜;i�QT˵@V�*��+��V�38����ɸs�m�rb��m�5:��+f��t�?��r��?��!��rB�+���N$&�G�/�E���"��%���e��(���l�+���4��Ԯ�t*/�6 +��LO3�-X��Re�U��x�[9\3���Ě�(����<��a�+��Ӎ��8�� ��$CSEx�ۆ.b��_��j�э!����A�TA­B��(��:��H�7�$�k9^����N�J�,
'�(�T�|��c��i$}w��i�X���7ƪ	a��E�3�w���l%�����s^����Ev*���0�J�`��Νᇵ�]8��\h.��4���hI��~}�X���3���m��?�#p�Zj=EIB&ai�`O�ʬ�6갃���r0�������Za��&?�

x��������[�y�	��&P	:W�E5��Ě�Q���m��+t͚y3p´pk�F�.�+�ޏ��h�y����>&�Eթx}t�~�M�s<�O�|�$�k���.L�*kK�?�[/��k%J��C�_��Ѥۀ�qA�g"%Ί�����ơd��y��j�F	��'���|4�e:tY��C[xޔ���?s���W��&�=p��w���oi���:��s�@��@2����S{Kbe]DW�{.��-�%4����U�׋��ڣ��-=H���=K����(+�\���5+9=᧪��NYY��Z�G���r��͔���JG��Z�"���k�$��uAK����G'N�����;�+{x������*��c�qz�\���	�鉂I���6��o}�=�����I�>F�9O#9*�#�	jD8�+?���-�bViDě��}�/�G��V��2@����mQ�aJ������.�e|T�����6�L1�c��M.V�oD�B�� ��k�P'a���=��a>�s������$!�����ОX��s��ΝLEH��ވ��2�f�r�׾�6�(����u���:��Z�����s�w�'�Ȱ��,�b��]��Q�f?~�tvGO�Sk'v?�5���'TF�s�j�F���n�A�,ϴK��h�y���-��˷X���6�4T�-	�������k�)ۢ��X��s4��$B�[�$t�����nQ�/ho�r����, �8`1A��
z� �f.̈́�H<j�i�T�ʂV�"2Y��lGȀ�#6�Z�)�� �2��c�~��N��n[�ь�P�tu����)����S�qdffԒ�#cp��<s3�X���y�D��7t	�4��.��|�ȍ��Fa�ό�Hw@��y����o���g~!������o#Jɦ�ga
��l��x�$�M�ȑ5�7GWx�L`���0ۉ=0b�v?H�6�r ���ژ��8��!��x��G��g��\E�?:�6�O&�����?�!`!���,�1���l��WqS����*FDǰ�C0�-Ӆ�T%���(����U/
p=��|!!��(&���h��޴O�l=��a�����|}D������#݇���t���2�.�,�k��g1�F?�P$�H���@�w�������c��R���V���H66������)���β���j��C&��;'޶S+g�H>�O�����]k���t�!�;�E|>����1�滴����X�Ő�{sJ+���ۣ{M�Uӱ�q�x*L��!P?���_4ۖ9�o1B����}�{�h_  T���}���󇹍
�+���ψ�ܢ��uT#A���	1���p9Qxqv�x��4^��O)��&��H����i���XE����8A<�Z)-�|�6J��	E������\�R�l���Kwթ�����.@��!>'m�$�����A�#�N~����PW�t�
?x!x޾�3;�Z�@��P��Ӎ��p����9gX�Rc���&H�B�3�W�֏GSS�i���i�.D��(01FA[�{���x�x>;��
�C���j����z��fGY��v���d�<�^��E��':�� �;�[�bc�"2��ެv��h�ɛ��>F�>s)k۩������ԟrr	��SpN��A��'�!�f(�vdr`��f��=���	ɗ�8,$M<�{�O��vaf��H���|.��1���c�V�y�+g#:����c]^9Nz�Jt1�Br�G����ܽ�H�9ڝm�� ��f���RY�S6,9��
��LRhT�^2W���@L;{:�����	��qTAT�yĨ+X J�˱����vh�l��=�%�ݜm�]��rA ��~A`%|R(��G7�3;#<X�@8w\XX�5��W���Kzݵ�R���|�;� n�4(�l�KVl�N?����-���p�������cQ]X�􀂐m�9=�`����E>��-�`��{����A.D�GJ�����5���V%/3aw��G��CM9x��҅��9G���	�vbN�FQRp!���^Z���R�u����}�ͫ�Uu�\��X�c|����J�QF�����~���k�V�19
��ϴ�iM��R���0�ed�c��db|�v�&�������F�C�#-idm�s���%�h���� �Ca������B'Q�)G}���GC}I�����R�NMaV���iֿP����v���e�N�$�Ü���>��bx_M�|y�g0��򳛀.g�!5�*DP����)��::�Gĸ��_lLX���	.`~�v�T6ĵ�JQ������i�y��YVMd�J2_u�m�up�I��n�ևS����!�̼��˵�y� ������0Q��ZzЛ4&"N����Bo�1�7���Ҁ�9��������$@�`Ћ�����fw����/�î��	�IƷ�%�S�.9C�D1���U=B*,�[��H�#�)��S�\!i�/�'�.)���9V)E�bg�7<&-�}�фte�l��"�227 �<#��,5'���^e.�.5Wl%dP ��F�0M�\���ޝb���Zhd����S͟�(ш��"Z	����Z��:���ݘ������rC����➯�!��M�st���{�G.�#a����N[.Pi�h-���[�<�< #p
i8��}����ρ ��qM�z�%U�jʰ��SJ����/��dҦr�?MCR�;��Rs��U�Z;9�� �r�x��R�|��KU<KZt�̷��`��r[/v�}FN������n���0�LG.
�2�켜�O�V�$��@���s��i�\#e	�P�lq�f5>�ߑ8Bd�bPKx�?�/���'�0`R�aF�v3P�M��V�����5���2��j��ֹ-!�8 .ܛ:ޜq���h��Q������M�A�1 ��w6�
���<8
������ǆ�ZS��Mִ��7�V�obpξ@�a�x��;�&f�D�S%�O�	_S\
���n�02���~͖pudf�[*�8dX{ģ�
�]/���_4��%����#�oM�%��l>�?�܃�T�B?+W�V�	d4��g������������Ʌ����G�J�z�S?~/fz�H4���{�}zXG��ܗ�g�z���H��B�US����v߁vcW��)-hВ�_���0��5+�����W{C̫^XmVL������5���O���euP[M���B��G��+o�"�J[�����7�_tҲ��¨Um��"8�`��Э�^3
HZ��h�X�5������ݿY�;��^(����ֿ���A�8�:?���`�����f���ɭ`�.�O�XC�Ѿ�>�/=#��C�l���^ ��s���$�l"F	Q��u�l�
	�TC�I$g��XFal��A���*�.O;֬�!�c�gu�^��E��&��Yo����Ǹ�+r(6ABY�܇N��i#�Y}"!az�&2;�G%�7#W��I��ӻ���G$s���������
!G�a�Mr�mKp'��+x�8�y��YjYZ{J����������9E�NV6
B���1]8�@��k�*=w���W�]>�����3t�jH��AO�'���>"*c��j!h�����S�h�NV��f�S��=u@��#ÐBk�谌W��frr_x��F�aLK�S��R�+�
�|m���L �rS��\j��^�/~��=�&k۞�3D��8������VC�;�i?���%a�,�_����-�g���&�ah{	!`F�NG�|�O�`�FR~�T�D`L�?��><�N��+]�k��jU鬼�ۅ`���t5��x�h[LLA�]G�X�\i�e� Ăr{�|:��q}(]B�}ǖ��B�MNh=ϙa����(���ti��Io��x� M�����4ލhg��aڲ�A�kwbS�F ���5�Ŝ=�z�a�DI+O����X$�a����g��;:����w�zm;Q���!�e*���1oRYS�����n�~��"�+�T�\׶����� ������̕����	�����v6�Z�̨;�dV���B_�5�&E�T+����v�y�#�P�G^��Rڥ�bt�%<萊�P�Ż���V�6<L�$+� �\�C�����d���h�<� ��<P�"�J.���ə����y��m�^�B���=�m����\�z+}�3u�(���nq\�O�0QaR� :5R�}�\Xj[�[}�cD�d�d4G`o��#��^Mg	�6��B���Q��H��eA�Lp�LzW��${n���ߛ�[+B�! }�Y~�0Q\���,���7���O&���%���~�t���$���t�`B�`��~�~�v/��k���ÒTǾK�\;�Q���p�Z%��.fC�
��}�clKfXz$8�[�:=ؙ��aF�c�W5��1��$���l�s��\I��"	i�V��KJ�Q"E���;Rw�����-��s"�'�xZ��7p�4G P���.A\� �.*�͋��QE�,mi�n�8�A�B����U�=0q�#���D��N��8�
*T���0��Ge����2�r-8pT&Q�J��W�"�}^�_SQ@�{ĻD����Wn\w������q��7湽�wp���?G��,]ثp?Z�wEC���*�*]��l,���釈&�yS�Q�2c 
N�1`Px�TӒ���4C�Z������_��	���	�yb������ҝ�0e|��:=��Q�"��R�:���H��n�4������X��0^��d��,�����!�m��3RF�0����D6�~�W�p L�+�֧&r�s�	�b����>]������Yq�t?�kq^��7��T>��M<,+Dѫm^��f���^������2��`�њ�Q�C#(;ھ�+c'˦�Oéڻ��fO۟�#m��R�0�����m,Z��^wA�l?C��L�P�� A�1/�yյ���2��Ƿ���6W"xo���x����r�zb	�AL�s>Z#u��4j�d�������'��3�Q�([1��ڄgk.-��c<(�)D�.�XP)����s�uW�\f�VM�l��}�}2hs��U��g\L��>���V�p���pW���cD �� u�lI� �D�JPʨ�iœ�D>��C����8�Ǣ�x1maB8}à�k������TK%�I���m���+|z�Z&�����-0z>�~N����w
����n�3s2�8/[��nhډ�B�ƽaX�"�ݒRB�VK��G_��a-i���)x��ӧ���O'��OSut?m�����LԈK~+�u����L����͈񱐍���?Al�K�P�Ti��R0��b�Ypȡ|H6���I����$VP������SD��L��]���#�ۛ���Hcʅ��]|�,���i���ҟ���@H�M�6�nBٜ�h��N����*�D���8���`�{�x���`�� ��d]	<�.��Ai\�up����V��P3m�KG�Td�{��f�p��HJ� ��D��$~����C�- rݝ�X�{d��ޔ����{�;��#�>�G͡Ǐ�����E������>\,8�q�m��� Ks�:←��]�6�G���p����M��
uyY �~��s�W�'���ְ�/T�إ2�b�i���ҧ�R��Ψ36�nd4��.<�F3���d�0摠pŌ`tDm���&YBȺܢ����_�z���X��� N��R��T7/"��eF{��.g��oi<WN��q#�*�%���O�tz��.�MY���>H��;;��Ŷ����HR�`��'�����]�
VÉ�i� �"=?wV���zQ�{����}�yB��cz�Zoq��s����mG�9�i��+��~+�ږ�[��OQe�P���Z�v
<����B�������Gqg�ʁO��}���I$�ݡ��q^����{��s#��~�jx�&�|"����a�/Ѓ���cS>
r��b.�M���KG���A���:��t�1��[6�X��φ㣤R+����e~N��ྍ�;E����!��$%!{��cD�]�F����k���S����uIX6�������;s@ly~uqc0�+�O,��[\�`���{`���,L�b*r�ζ���x��M\~�GQ���߲A'&$��ɴPonB��P���a�n��\�{k.��|��O��=��C����OP�Vy����~�3� {Q��v�
�Z������q�s�s�S`�UNv<����*�����neK#kgVI��s*�s`�zR��;`!��E��xW�a:r�?�8�]έ3s��^cGy^{) �GB�����V<:m)�M�j�	0�s�ӧ�[(ڄ��:y�c:�3fS��!�� I�.�����Ip8�9?7j4R�'i�:�͍�������y� � z�����`"�v��T\_� ��mf��b�ը�L�`�B�3STo�S"ZMw�,L8x��c���͛`�yy�##�N��%�f���HFG�yKk7Q��� �Ԙ�m�'����4��6@s���kfp-�r��79�B�hb6����xP��.�2l�*�J Cp!;��i�!��Z%F�C�"��~��&�W!77 c#w�5E�ejw �d+�b�H��Ϋ�H�����������6OcM�`�	?yd��`�-�|�ؿ��8N��^9��!�H�	�N|�ՇW߲%F~�mwm!i�~}$�Н�]��E�XB՞1'�>�y4Dh��[Mp����)��/�l6�f��$��*�*�x?r`���� ���(Z�ɜ�̅_�J���S��in&��:Z�&���ke�� ob�,ɇ��>����@ �� <k����%Q̬z_��sKf��Q��7�+�J̟�U꯬�/� o�}*����!�|E����C��LZ�}U�u���FI�'��]b����k��rh;ZpX�>�n���� ����o�,��1Z�=X(�;���5��\�H�7��B��F��H{�p���m2�ܽ�v�
շ3m:��^Z��	����g���Q���>���'A��8�*�����ˬ����X��K>�%�[�Pk���3�T�L��'W{�i��7jY��ol<]��H�hHQ��G�D������­6rK��鎋u�e�@�/ݪ�2��"��Uxm+;@�2�U%Vj�~؅�c���9�&Dk?�]F���6���+�/�x, ���*��w��6˼/n'�w�@�q�� �
��\�H9ȃ����|�f�����E�7`�U�����>^>��u���3��I��*��x��Y�z��+8�_���y|���_����8�}�Ko��� #�1Q��N?�HH�M/$�L�f���Ј�	k�+��ȸ&��h�n͗je��s`�|��)�$���j/���������yl�x��^DρJ����t|ز��W6�zO�~hc,�5��X:7�4����'���&�l䀝`�j�v����ZL�cN�ڡT\�_w���9��G*����(�9P�\��pY$�����-�X��'s�i,W":-���mZ�aG{J�KmTghͲ��}�HW��zҰ|q����Tne��Pg�)���� P�7h/��,ob_~k� *�lj�-Wh�����4�D��Vx�S�j(��db�]@�]�
���||M���z�/��F��y�^@e�|\�N�d�$���i�r��cR��ݐ�P�wd2���6�=�4�v�jk߱��e�k8#^�Lu{)���S�"�k��j~x��u,S}i����Z�;��i @����èY.y4��,Yl�ݟY�V�i�չnj��%| s~���R��㣅��,�{�b2��.<�n�<+Q��g�f�0D�O`����+�Y7%����a�������P����V͔����66�#0��YX���  ~6|� �����d�:w0�v��*��CiҴ��2i����OI	m��etO�}S����&�u��L3 ��]��nU˗��M`@ˁ����z�#b�B<��H��E=)A7��j�DvQ� o��6�����xp�{z��^w�.W��Z<�l��P��1��$X���!'��It��7$��]ܜ�1�]L�t@����LqT� >v�J�:�)�DǇ?Ѥw��|�q�W�,�����(�@^��j�Q�V�whj�|?ӟ���~&?KZ���7!�H?D����&�)ѕ��f�2��4
q�i]��\�M��r�J�(���kD�	 �EG��Ⱦ
!I���U+2���!P^�n1��)A�1�c`������5���X$���&������S��@�Lf�k���P�G��G���5P��d�E�Cv�D���Ʉ�d0��:������Y�&���;甛�vjS��*�S�C��J-�0��G�½�.'�%׶>�A�1�@a��;�KJX$�yj,k}�y���f�x���O�,�cωn�[�}S9��DɅ�rD�^����ڝ���u�z蘒eҢ4��֯b(*�k��="4���lӣ l�At-�ϭa�#r�%��JY�W�yc�<\��M8�'�c0q��I��t��璝��N-15D�V���Q��S.��Q	E�)Z�)�h#�Ό!�`��r��ǘTS�����z�����Vo8�ei��S�B��@߽��
���|��Ji���Ĭ�eT-i��+�i��Zd�"��MRM(z���U�&]eW騾`���5�`N���=ƝAq�S�:bbd��x���gܳ��kp9&=�K����]0��L�����lh�%Iu���sR |(0��[�����@)�u�$F�Cp���;�y�����eb��1[��8�dN��+H��3-�������~�����KzK�W�Y�
E��o- Ǒ���I���Y���X_�J]�t�4i�o2{I!,J�୻�����r����-_��>���D�c��B@b7a9:���C9]��kM�x�����r�yR�A��x�P;Q����W��h���Yx�l8s�/���7���g��BD�м@o8t�},��	�� }����l�N�JIk�Fa�B��=��i,s��*?��}�_,�N����q(�9����d��Oh�"�������}S�c *'ed3���w�\�a���6�Ql3�,�����9B�lǷ}ݚ�H#.m灕+`��x���Ùf����^|{o4�b�>�{m� �q��V{(9��[醣�0Z�>�����qwB�m-@YH�� gaF�⢲�T�v
6fa��_�447sd�I�����Rځ*엛�#;aa�.$�'X$��aI4�!�R
��:��?*ݐҌ�]�6{P�u���x���B���������I�s�.c�Yk&��>�'%�RE�F?̕M\��?00�L,��FNr�z6�7�l�umW����1����V'@�ujA�
��4o��H�w�NM�l$+T{ �T.�7��:��|�M$ˌ��#�֭h<4L6�$�A���
%l�a%��̇�+�ҳ\��f%��+�咞��KCN݈��Ur�a�F�;m�<��B2m@D���j(�����O�G�IA���2��ab7<��|6�=��q�k��W���X�%�� .FUMV<#��Q���8�V
ޔ���/��:�6�Y^Gu��0���fA)���������٬��5k�Qb�Zd�wo_�K)P�C�CU�Z.���?� ��}5D�����/ޒ����䍻E�������%0�6ʑ�.�)�*�JC�0|p���_�k<V��u6��@l5�u��e���Qg�$�������JLmƮGΤ8i�h�֖5�_�ȞXX2���G�ՙO'�M.����,Bɟ�F��k�q�>�R���1YQ���٠ =��m:Xn,��y"J�N�Ŧ_Դ>>�8���l�Yʂl���o�.�#�m-��8�_f�w+�W�a��Q#�rt
@u��f֑�� �`�|YD�`M����˦<u���4A��IEn pH[6�^�)��>;G�+8�r�;���z�T����*��a����;Vl/ـ��H�Q���C-hO�����Vx����˂����4�%�c֎��@̞�j-(�[�X}�����'�e�V!���A"�Cث���=ϖ
X,�G8�m(w�1��f| =ʕ�ʿ*t��>7~��搘hq�{�$;�]��4�q��^EK+b�ģq`�K���:x���=|}��Ѫ�F��g����*��K~n����v����hH�}�8�D�X�F�d5�)$`�����N���%Ov�׊a���� �9L��M`E��h�P��]\@����7��m���C�K� gˇ6���#�GΞ���w�Yp(��ȉ�>�����1A�;Z��:�ѓ��n�߁=�QKW���z��{�~ͺgaJEА�F���po�CnJ�V�5�FP���c{ܳ8��kr��XSt��޳�ir���Ń�dZK�]�w�`G���:�������G&=,O�\�{��E*�$����Mv�e���C�������bⰶ�vl%���L~:O�A�e!������[�r�-'Vt>���{��7c�q��^>*s�����{�r�w�3�au��t��8��Y�5[d�p�t0�ũ��-�-��O�b�WNT e��Ju�E��(�H���Gr����ݵs��Y+S���I>Kb�#�4	j�3�n�w�g�إS���CԽs�OvXq9\آF�3�Bn�/�&bl(��7;�iN�C�@��������.��O��^ }E�v���B%�uތ�{4��� P$V�K���:���mR����x;~�Z����t�ر��a�>.��6e	�qb��3*�7��w��3�2+��?������ӥ"�������U�hC�\�S.<�{��^�
@R)W�(�
d��Z�GD�t|�:����	�W���a|^����eF�_�\�x���S4�7Jt/��o�c�ְÕ�ɸ���m[�u��Ɠ�>_1h��R��H���k2��v<'���{Bp\�^r��))��o����������ڻ��+�dK�%�=P��W^CV���ǩo�p�b��hh�uT��v�
��OL��=O�c����Й2���3R��kl��k�;�� �9���K�/�IKB��GI�����	��|�����vN8��7���
��cj��Mq��좲���i����,��=]=�_Z%���
c�a�щ���/��a�K��(��SsNbSl(	'ݨ�!a�y�}��!��H	N����a�F'5����t(z�p ���T#(j��p�Vt�֣sӅ��;��r��*��sRۘ�r2�j	P�{��r�!��nl�`fRQ������d�׻���F��C�㣪ˁq͐t����O�3�����]df-k)cx�"Ѯ=�J��B5��D"`H�_y�������є�> �J�[�	�� �7�*�E�H��Hܪ%�Y��e�_}�i���ĵ�@"�Z#k�,Ƅ|�/�.���nӓ� ���?�DD��{�a9^��`�pu�s�i���bE�y��B��H�9|"G*]aOa�$�>b��e��a�S���"�_�3��Qi_�v�Y��`���+!�Kg�sC&����V�K(i�x���l�>dϸ�.Wa�<���^q ���{V� �bɧd]e�M�DĠ{��r��u����{+f��RD%�s#Հ
wP%U�X����J�[�}?5���c��r���d]�7hI�ԗn�x0�G˦��⚾ѹ��:?�u���w]��YW8���'�,T`q��=�"U҆zh$V~�L=�+�ڿ/���KVs�%zIO\���}oT�9aF(��6��o,��ķ'NI=8a���O�#A��!�BHY��&�hJK�eE�9E�����̑���>��H�{+�F�� �L����&�ػ��Jr�z���."��g`)��4��a��K����C��}?��Z��c�Ia�J�Z��M�͘>óU�D�*P�}�v��%:�)��o).������Gx)��/��_�1F�9	`DTlҞ"�c���� ���0����j��"pO�,�v`�r�`�p���Y`ڣ��Uc7zt���"RK�;�ԯ0&^"�m͛ n̎��X;���xʈK�w�O�bt�T;�u�Η�3�3��_�8�l�T�q�*�B��f��a��@���9ok7]5Ms�H���y���߽&b��Y�h(��N��\���?�$Ŭ��86���7�?�$���0*�K���-��g��v���,�Y"�������$`O8���~J͋�8�Ǻ��+�l��*3�$��;�hN>�ҁU+�q�!>���327��EɌ�nc^rO�]�	7r�]y66�	�dӰ���Mr�+�`zϯ=7=b�d�U=Wy�G��a���1��p�>�v��ժ�0O�AubȪ�{4��}�cylq
`�	'��Kd��tJ�lϣ��v!��,�Qx`�yyF	[>�r0�Nq���ߦ��zw&��⽷�
�|5Ta�����f#�:��H��X8D6�P�WU��L��OX��V:\���1u+�,�يߤ�M��I%�#Ѽ�#�<+;5Nk�S�+�P�'s���{7�AY�nY�ԇ8���|�P����c�����]ouX�#�%_�W�-���#X�	`����o�D�Z�����OU�-v%����n��F��=��2�ǃ��U�ݘ�J��F}�Į��Ĵ.�+�dNl�.#���N�:}�!���� C��ڪ�3����t�xo�0�,�b��-c�k�7o�A^ܸ5+�G:x@��/w���g�w�`8_�r�1�U~�k���j���x�K��~���x�����⮍\�KM��7���z㭓Q��^�^�rL���p�9���o$�!�mRS�;��@��8T
FĿ�0�Y>ve�("!�1[9)��n��K���=a�z{���O[U�ц (xd�ѩA%&u�Hw.Baa0C��$.�_�(��� ]j.�^ЭQ�M������b���q����ɾ�5Hm���8,�������a�%a�����+ �;�rK�>w��C������ō�H�p�u�w�2�����e\0R߹����á=r�����yq�BDj< ���/��n�m���c�b��L�Ӑdxs�[,�Nhzu}h(�,�A��j�i����$F�%�o�G�һ���kGM�W����+��ݽ;�������DE�u {I�q5���P9�t�jg]-��q�vʭ7T��c��Ջ���LkÆ�>�ă�X>��5�p�c�\����+�X�],bq��軝 �@�!Y$vΆ,�:��W��K�lν�̅?\Ò�TAb`�ld��^-��#� X��Uٓ U�+�G�I~ ��q��iӹ7�[R�\?w��{!1K�"{d���"uGo�M������U�mϙ;]�%�R�Y�X�?y���}��� ��.8Nƚ~K�q gʉe}�$��gh-Pw�����Ck��Jym$
�<JW�F+��MǨ(�K&i�6ύ���D,��rf�#|X�!A·/ ��am6�\�6����{<~"��[�+´ �inz�|m��Wi�*x?���%�o�9� ��:���?_% O$���5ҟ�r�d݉�Sw!�%7Ne�X�p��p���(���Qi�I(��ΘG�S���!���D��������j�Wۯ3#�UiK�����<]�ӧS;
Kt������֊b 0�^.u����E�uш3�uOG��y�	C8�Pӷna��k�� 0�v���"���_$�DN�l�yT�����=�@��St�f$е�?��O�30�P����S���(Y�J�W-�z���&�#}�ܟ؅�(�7� i�J�됽L�7c}�r^�GZ�h�Hs���^��a���Aɟ�y��� X��63�B�W��h�3��U�EP�F�h��,.�_��=L&�s �[K�6a�p��"���褾pho�W��Z��? ���io����D'�N�O�+Y��Iw����o����ۀ(��=3�&��d�Xd5;���i|-|�
�f�#�j���ҫ�O�,Svyx�d��=�R�9�d��[��4�2J�W��5Y�ȯ���Q�U����҇>�h�!��H(��m*�5�d��P�_w���o		��d�*�N����=��T�b\��~���N�m����ԝFiu�:��]�O�m\!ƂD����h�^F<��&#��}cy;P���U��ì]��{�A�����%1��ro줞9�?=��}mb?���qeM�bA�W/s���ըx��TS��G-9G͗d�rڞ�<OW| �N;�Y�	wf���C�����Zd`Ӎ4RdS���c���ͦ���ړ��j3������w��l�l�>7���~��;�ҖA{� [hg��E!�˴|�v��sI7S��}�`L`��Őb�&:�%B��t�7H{��'�+o��� ё�T��}]='Q� ��O�+	�.��W���nx�-A�J<;ٺ���ֱH.�s�ɻ���*�@�@'wG��w܏�',��ې����&���倀���6힍`by�P���ڹZ����,����:F`�������,���Z�EA,v�N\��FN{��+��V�w�Ӂ�	X2/;���5ar;�C�K�*�S��9H�'�0 �U�+A8��Z=�U�i>�e|�ܹíX����q"9\�YDe�6{cJ���� �8��&1K��Հ3o��8��,��xM7�1؞m=�.�C����� t�y 9S}���`�}��K�~�B05���T9>,[TP����@X�����<b��3�]�NAc�3��)7�����x�>2x�wVVc}�%�A }�4F8gJ8�*P |��~2P��Aݣ?��^��?���`�pr|A�zN4��G��H�zAe�k(t�Ѳ�Oe[��n3u�+�j�EF���G��j�����S�������C�.b�t]<�Ye�RDf֎֟a:�zX*�Cs}�]EI�V H��ȓ��巈q)A<V[·ęhpK�i�b��|`��5�^wS��g�v(��4N��������.�s0S@rh�+�_<��&I��	��Rc �������?�g�1C����s<�7���v=D�nb��Y� �9t]�ujy�ÄmA�t]��t����D��Ws���M�+XE���o�F����--L�>��ɹ����Y�t�7t�%݂�(�I�^�P0C�h\M�0��6�3�e�[;G�Ǒ��X�j0���~�	���8@�Ȁ�,���qW��5�pu�(�ײĿ[4�A��HcLb��坉��k�&�WY�Q�V��_+�0ϟB�ڮ�"�?��7	�<��`F8�Xg�C ���7�rC����i��?GQ@d�JQR?�7���͜��f5���ʶ&|�B����c$e�2UB�j�8W�>]V�c�b�{y�-ci��kVd3��H��ʟ��p�QpU޹�]��y+>�)m�����#����R��hR��z�-��Pi���[0fTA=��Lw���q�ǎ�A����P��J��t:<�d71������Z���	 P�����}&�8���8�4
��	~œ���i�)�?z!�
�5� ��X����t���*� \��T�����v�Y��/VX����_��vO[L<�A�fm:��qv����)�d3�����	�nA�"�L;7ӑ���؋�A ����\�53�� $��[�V�"~qb��S}H����W��c����sU�4����/���T��M�`|��M!K),3 )�8�M/
G�ԋ����m���l�c���k��;`�}tP�J�}�c/�?9-xn�F"�c�˔��kI��K���3��$ڀ�bY�>�C� n��R��T?Qw�G��������0�g��ҏJ���Kc��h�*6a�Ը�3|au�,%z��vHW]���/˿eaG��qe����ʎ�����M�(��wƤa�sƀ/���>��zjwW\�t��٣q9|Fp3GA����5�� �b(iU2�XEp'�������B^ƼqUC���{��
{x=o�u{�OF�q��&�d��<ӫ'a�H���\����1�;���|�q����:���].1ގ-�بs%�$@�i�V�y�.�q銭d_�l��2/vQ�}Z��xA?E�=�}� �;�u'-��_x����2`at%"o����t�'6$���ں
z�6X3#�_�z,�r��O���$hV[N�̽��-NU��S˦㢶SG��@U�UD
x-� t����/��� N9e��#K��w��,�P|Fk?���\U5�8�d����P�ml��(��2ղ��%!%?Zu+���6�J�]+2==�\gPY�	ͩ�C�.I��X:�ޭi�K�i����g|�D�B����aB���#I���I���,���R1ĬC<��B-�ߎ�紡VH��Ū
nFJ��P�E71�Tm(*�����ˉĳ�cL8&.9W�R���9S	�8�@�Dc����"Bo{M|�[)�;x%m��M��]�4�P��@f6->�y�p���k���Z/��; �H!uXAQ%������W]5�Ym������k�Xs�
5�[6��j����D�p��t�A;��g������ �F`���3s�j|��Ŋ��n�";ˬ�Q�{i�Ø�HDq�&�*ăc�ĹYp�Axh0�n����/c��]ܨ�E5�&�/%aP�( q���f�uEݳSA.���qlb+��m<����jboܿ���q�2�E@Ơ��(��S{��E��=L;ۓ5Wpwg�5�'H�#���@c�/�%)�3�� �D����`V��m�[����F�(D����$���fP�A��,�c�Q%���Z6 F��s�7rN�ˑ�+on��s�^7�pzeAU������^c����66����x��m5��0�K��<��t>���l�zZ�=��BU ^�{���a*��X�֧��/%M��0�K��EEfL���LA *�~a�R�ltԚ<�x���h���z�3�mq��$B�|�ǬZ/:�һ��D��}���4�Ⱦ8��w��j͗ Vs�Z�7*ܮJ4T�FR'Sl���9�e^��T���pJ��U�>l����@2�A�¿[.�<���4}P�s�&N���+p�!S��]8�"�sY�X�b.�'"o��&���<�D��D���=o���:�*�e~g����z@��F�cf�ok�_�H��S���:05$�9(;WU8W��7D��y�\��Q�w��i�(NC5�Uu�x/���p&&�t_����cOeG(9���r�11��yM���3ա�6r1�$=>��K���,we��%DL��Y!�Og�5���@�!g�A���W���#�I:P��Yy�O�����Ϲ���i��ͬ5�?;���{�s���>f>������c6��n�;<�	4~ޟ���d�~�kޛ��D�T�rZv���f�s@-^�Wۘ)����Z�c��n�H1Mo|����}	� '6KV@�&�+}5� �c����^�xG�H`��k�%��!�:0N@����*����G�r�(���BNsKw�q������C�ȱV��.�T"J�H�$ ���Z���q�Tܽ@����W�����#�0����魪�אLO������/�Y�~��u�����V��*�����+U�F�]�b���"�ua��:0��q<��%l����Ϙ<�so�o/7iC^�-�לΗ�$IQ%���Mb��D���GUP�\y�x}�_j���F8��eT�Ri8i����%��L3�������^�Vs	N����d���*`(�{�n��d��zl����1�Q����"��rs�4�d����kO�rsl���և���G�=���O;�R�5��튀��j:���UB�K�z�ϢP\��#��
���,�sA{X��;�����\����`�6V�e��n_������y4F�˧�l���=����:��ͫ�־�2���7Ό*�ͭ�
�,0�,rI��*ǰ�lfyb$�ԯ�@�U?dd��^tC�o-��
�1��5���%`����3ٳ9�*,r����jϡ���`����+���Z&���H�7VDg�ҊK�t�����:���{��ض=}7���B�ܦK�5��e�u����������*���F#��B��Lz@;�c
����J~b�Q�8!6����BW��(�̌=j|e)���h(�f*��cP�רFC�����Rl�Ǔ�s0�y����O�.7�'�������4�r��oi<`��1�)�q��
�%�L>?���Y�e=�O�5��'��<i�N+�=w��/J�{51x"�L �p�ŏ�I|ס"F2J�\�Ӡx1���7iM����h$;0�x 캍��/gELe�����g�C����V�N�~A	I�[g[l����I�����̦r�Ur�@]�L͈ڛQ�O�zw���{���)�Q9-?qƳǕ��kd.-2U 0Cm������*�D��x|t��?��~M֔mȘī��e8�Ō�ϡ"G�������4y��5q1�~=1~?}�
�����b���"�".�{��lx�"^d7�rk$�S��Y��P:Ã�����f�X�����`O�>x��!�. +�݄�ҲVGv1(��}V��(�{:�4Y3^�_PI�� �:)]��g���u���⽼�1��e/�B4b��9󎵖�U;gd[M����,u�.��|Z`@���c2�R6�bЈBJӨ����l����c̭�eқ}����/�)_t���9�4�+kLvn���2�:bt�R�������v� ��!��sr�/����&�� I.��3F����{O;�8�<s��؝Z�	�2�:��tjj;x}d���ݣ@�P��VM�a *�.>?w�e�"����э�eʞ0UYV:~DoƁA��Jd\ZM��h�O&��
�'�^���g>__;s�$�8��?Vȧl"�}�!��I�d�Ã.Χ����A�pxn���z.Jo��׼�P��0���o /\[��;ţ��n���%��w���H���Ø����델R�����@�� R�BP�7@�8��&�̅�i ܢ���o|����G��/�2N]�]X9���6_��9�%{How��Iv���P�V�>3�z��k�o�~R�o�S
^����ȸ������k��v��LL������7� �q�3zN��hza���
�ǑĶ���&5�t��N����	: �����Lf�_���/�K @u�q�n�2En��tM��7f	oc>G�7� �[GD#¥w���S�+w���z�R�/�j��)`�k��T����XE7���!�֮�In�ٽu���7!� ^�g=��,�b���qi���Eh]64��������`<��s��	�J-L����̤,j�ލ��و=����"�Ά,��BǬW*��,����M��^n��> �t)���}?9.>_�# ��ѿB��bm^\�߇�!���/ME�/�����w��X��=�ᱜ��9(�� ���D�V��ʮ�Ar��P�$�!�/��h��Kk81�D���m��=C�������][V�t�F�yh$B3���U����ـ2l��7x%�S�s�g�ʬT5��][�����?y��r.�؟�+#�R��I�+�"I+���+��&WGK�����/��0ʻV������q	��K�O�N �P3D|A'��\�z6a	���*�+t�\��MWe�x���@�Ze�qӔ}��`�}x���;��r�&�m�Q��W?��1I�뺡�",�L�䬅O�J-T�9jӣ�]�1ՎX�AiC{C�����;��J���,y�t̚�.�+����t��H�i��`�"{f��:�Ƴ���cl� V֔��S�*��g�c�Jeg5�ew=6�#/�W����.dn�|'��IܤI�d�\�<�q%�K2*[W����$��6j��glm��|�7d����2>�&鮨;��0)�E>�H�ݸhٶ��PIj7�o޵�d�D`��� v��TY8u�}��3����wu��c>+%k�sv�l������Q W��-t<i��WJ�ޮ��<�Ak9S&i,v�AK�<Z�-'Ws�-���|`ލfZu����
��\pL7���5�{L^l�mV�n-Og/�rz���[s�� M��1m¾y��)i���{t3�E4מr3''#} M`um����/��iD�U
��h���'�'1fHf�z��_�vE[���a����8� ���D��[��r�����j�avL���x3��(�^����W��ĘnW�a���c��������<�T�QD�vr0���b"ϻ�A���w�P�T����2���=� ��"E��d�a �T a{�~���{�h�� �\#=�ݘ��[��.=?fnԶ���cX��S����hHv���Dt�������_X�8A��a��*Ǌ�N��ƈZ�T�Va�/g��B��?���
�,�A�3R�9}��>K��Ʋv���}@�7K�v/�X���{�j|0ڿ0�N�׭+�+�^�f�4.ǘQ�䐨�Tt�5K 5����_Bq�~9R�׺좲.�!8}.�U�u(!���b������Z
N�p���DsO�����J՝4 �V�����(� <�RKs���c�9�@2ܖꎘ0C"��4^k�ZF����3˅Y��C.�S��ޥnn���o��ֻj���=�C`��c��g>������T��4XUXj5G[�H�w�W2X�w���a�h�&4L�K}VOJ��A�% ��C�K �q�d����o�Fj��׊�IŌ����������������'�>y�����k�ሹ�c���T�W��X��B�����45"[��]�i�竝��u]L��������I���9��p�;q�?��w5ZX6�|T
�'O�܎�#G�2���[����2��Y��c�Xi�ܳ�c�T$�T�{ �Ks��������xKZm��!O�j�S��,X��P�P?ì�M�>�'.h[�->r��G�k°���C!�!4K/�$���b��g�`���Z�m!��T�$�H.53� ��O��I��X�(ëfO�=+Y�9�1���&�� ���f�`�'��:mn�k`�E��fn�l���gzWI��k�������P�-��[�K�nD�0�>��]C�r;[�+���#ҥ40qcqqN�7 �cU���@ʮ7�i�����b���4f���6!��r���/�7"=?f�*;��-T�E�>:��i�`t�׉�Z��@�M��o��I��R���0zUW�n�w�їBȄ��I��
/+��A��{�Hw�����E뢣����2cq�e�5��y�5N���e�s?���o����0��KZ����`��o��`��WOK(��ϳ'%�L���=�E�'�b-�Y�f�y��A�?i's2�2Ř�4�80/3���\а���2Zk�s�������Ԇ���$wq�40�^�]H`c�l�!�g��X�p��zz&���ka��Cn�k��BE<��t;���h+��j)���R*���Q�o��M��:���NܼO��A3�ϝ�J��6���o����֞��l
�~�P���!���Ç~�c�4[�j�`���� �`�@9��Dj�@��&�4�ڢ?�\`B�׆/<����pl6S魊�����/�{�w�#lX��ǀ��/�]��3���+/st	�np�<C���9���USF	���;Q��>+E%���j��q:}3B���`\�bףC_V ���
+V�SX��t�I!$Hb��"3��o���G�y�-���������td@!����6��&��=�=WX�a��r>ѿ�����D΢�j��(���o �$��a$;¸Q$%의���(uZ^�2�p����#�;�u��G�������|���`y8fuy�%ЄDאR�Ԛ������1'�Q\�<]UT~z��+#���@�M�I-���C��C�v�� ��$ջ�����d����1A�`*ܿ����F���qK)�?1��0�䌀lOY$~o�����'�M��L,��~��2�Q�����c�I�m�[<:G���w�N��6*f��&�
���>�8�(�8�"S��UQF��`;ڡ�>�v��hA#�UBK�G������o@@tL�puұ)�R
�B��D��#�Oރ�ȣ(P,t��᱀�b��$}��EҞg�ڕ��F$C��B���Ig���~r	WJ:�[N��]J.\~�vyx�5a&�C�
_�f�M�@���xZ�{$�&���,��Q��k<��B"0�t��Ę���R��z�':B��Nb�]=dr��V�B#�\cl&�co.����p�q������~h�Z�ɾ}s&�4!gG����1:�7�&2�ѥ{<�����8:Iw,vnfC��[wPR��1Y��^�ٮt��6"T�1��J��;���/���^ 0�\O�N����6>��M�Dz]S�<����$l�k��+�1��3�p�6�|����zp����� ��8O�![6�#ChP�^O�U1�����GZ�+�����㹃��`�}�v����Z�e�{1��0D�=�!�!	�$��Q{�qU�(��QJ�w���pK�d�7x3R�'‼I��U� Ҳ�b�e�6��*Q�rq`�H��BBq�Mfܩi}I���+���a��],D5�����Q݁����,�eN��Hx�r��+(�����LV��zEB�u��_����ZL��Lօ'u���� t�au��b�xv�w�7���roW�5�XYj�96�! ��U�&C"4��Ra���h�k��'Y�W���?~aUͳ�'>�ܒ���Ϝ7'���Ty4�v�<���!���]0(��AV�|�|>#�)�[>����d(S~�=&�.5�J�繚�x�c��D�Zuz�h\$ŕ��σ��G�)�Z�3�nrOu]�b��l5
�	j ���Tu�S��'�y�$8�-'�'L>���d.�IU�(�}�Q���(}x�2W�3U]��	��h��p�0�9�$����w�#���b��m;`�xa��[�>�N-0�-;j�\����8!o�pGWN{�%�\�4=���%6�Nn�u��^r�|ֿ��2�2^��Ǵ��!s6�`|.��E��}U�����N�c?D�[<̲n� �^�^�򺹒|r�dzpQ�:���X2����9brc�LdR2����\��Fig�_�}���i�1$��%��)������y]b5ʞxEI.R"���cy)1�a�Ű^HBv�<X���w�ɭ>��:ⳮȼ�@���L�5J�TԈS���S(J�U7X��
-���k�_��tM����/�a�����@���0��p�־oc%Y���Q]0��G%�ˇ����q�g��8_Zk��8=nwh��o�C��ϷC��
.��"�t��a� �~���u\ܴ6�y7xt
��0f?��!���������|�V�B)��ah%�:	=+b$N�;)���3����:�0;�=���쬒yszʷ�.��A����"��C>o�p.Y����n�����6����n6�$	w�+���^�\�bZ���`n%C1��I��(Շ���A�G&���t!��~H՞t_�"~4�pL&;eF�ö��J^�!�7,�؝���@���i;O�r�!Q�?}c����/+�tF3I�Z�^`��~�/i��U��Dg�m�,��*��N.n������݊U��r}]�	[��u�J�~�0������OQ����%^���+�2pŇh^|����%\G%���䥋��?�)�ۇN��� 7�%yγ�4�����!�w4�(<���]�b~]8(��������Ro�/�Ş�4sȯl�e	���#�qV�.9J�R�����Mb(���h���+A���C4$r� 7�c�,@{�"��.�T��I���]H�1EO!սT5������`yϡƍ��L�f����.H4I�=�4M��^�C�%��(��s��n�$p���x�� �/}W��U������P��d������d�2�Z$�2�^�P93�.��vR��½;Hc��O��H�7e�>T81��������uV1�=l$���>�1-
�v�&ya���|vg�_�?_,uW����Uv�o!GM[߮b{cĮ$����0K�z����/o����f����!�n�|���^��F�����l#����o�Ƽzy&% �f�Z��M�>.7�s;z��s��VS�f9�B}Iw,���u3󫝈�~R-cT��kP�>5� �4]�JfV���D�_�x#���?Ƅ���*~�(}7+�q�ay3��B�僯��b���8����g�+f�Tɪ��,7�4_M�i#|4�r(g�,�@�pT�%����W��OEӞ�Lkn�y>�7޼���Q�p�h����<��Ԁ����sӴ��UGn�S��8��Ed��	�V ��S�@��z�Uw����鎶�d~sW�.�-�iC�|��أFX�ZYِ��u��Q �y�b%Kk��a�(�}^�fQ��P�qcE�;_�� ��9������ě�����n5s"�<NG`�����t	�ԯ��� �E&s	��4=%m+�E�sp��j?�J��8�,��S��֍���b�h�eZ���D��`T�i""-�b+���x��~�U�0�z�;.��1pvl�2��X�.��Y�w==/IA���Qڿ��n���+�&����{4iJ,/��A�v��d\{�F=fS���I�7�,�\�!�k@P������|�wۆ6����ӗ>o�,��Ϳc
�~�jJ�m��K�?F�������TQV�O�KTG.�I�_�4�'ÝW�%��sc�N�o��U
Cc�\�����>�XR�TR� (�{ؿG��<ՄV5d�������a�;2.�Y�/�4�4Ϭ쎰`��r�8O�|u�S�/�1�$�>EW�Ů�Q�	FU���(�z�4p�#�M:?=ޔlkCU$@����袱-�v.�
`�-�h���0�Z��"Kw������.��Q�h7-� IT�%�{�=!�v1yUf�����n�R+ϣH6 Ԇ�R�g��*2�e1�e�b/�c�2��g��FU65�����1��G��:/��d<Ib�+�g͉�-�%VH: ���?hWaΡ�OP��3~Ke�|Ȥ�'È	�/���hJ��_^ϟ�>�!���o9�%:�ã'rt��}=��3�#���Zh��q�; ��]�\����q�q�+�����UY�W��ꐥ��I��.Z��ҏ@�:�_C��0J��x{9���(JO$��1Ԅ6 ���e��
j���7L�Q8�x)u��vA��Vk�F�̔������aB�Э���ܛ�����3� ��m+�PN�e}h��+�Í�iP���F0�gfk���'�K$`����]+���^��C|�u�F��6��ˊ���Zy���\��p7���ő���c�~�kX��{���Ȝ�m
31��!�|�,��|�R�;���#��V2��= ~D��`m�f�qĉ�h�ƽ�E�~�Q���-,ˢ�!���D>�q1hM�f<�1}������������� ��5_��0N�IмRwp������F�`O+��U6���U�0Ff�;�1^se�) С�� [�˃����M�~���r�~��S$P8G�%x?���/]�8V���9�^}�䲴6���xȗ>m� �(�p
s�T��,�0p';Ey� ����"J�uD���>v�h.){(���j�Q���������W�|�!��d��G�|i֏�� �CO�_�)F��ڕ����>}m��8�a� Rs�$�'"��町e�c��F�����Bv�m�r�=�M*�4XRB4hB�<0�P��0��r�˰��T��\0��/���
����)�_)ü��($r's�i� �A���:H��:�����mv�%��ڏo�����0vt���G/�-Dd�%i��v(�_a��j���jt���ؿZ����&\n�D���-1m��p\��DDeY� 0x¾��lǂr�x >x�bF�o����,2��@혤A�ٓB�+��ՈX�U��"30;h�j�hiǍ3\D%�jY���+IhEO��̗�X��yo�c�7�6��r,�����Q�OcEZ���e��cT�>�zW��QZL]l�6:��'[�������h#|A�t����OR��t��+�-2X��x�c�AlQ�^��%���D�s�f�&7V�fqYt*g�INd3��}}G����j����dm ^J{����Za�:��a�>�B��v�%x4@Ӈ�!��e������|�I7In�T�Z ^×��l0��y:(J<��+�Սm&���_dEe����8��1¥BP�\RL��67?����g���������~�>�9a#fxlF��/���H~F��8�)���yZH~p[�S9�v��H˗\�W�3�q��q�C��ˌ}�����O�����<����=r9��D�}����p�j�z�c��Fү����g�]���
V���iҲ��?g��݈~:�)��>��P8<�O2�����G�UW��������^�]7������^���k�=�u��e_�Z-�6L�(:!�f,��A�3���?�NB�|�>|�$��s�8�9����E7�t���GG0��!���"^�Dd��UH�(��7��ɏV�}��&���6��\[kwq�A/x���j�O75� /�b���m���c�N0�{ȝ�L�+�Y[�Q�ʠIV�;ޥWL;+����u����Y՜Z�ҋ�ɕz��M��F���!��~�c�G��w���z+� %&,IH֒��"�d���`D	h��!c��\�;;Z��Ӱ���#1�^�k�
�sJV���[� �>י�:b�&�<��6?����k�iF������� �BX�{\��Q���vt��)`�؇�R4J���� �5�kd���\�ϓZ�42�������p�%o >�a3�^O����'N��FE��}yb||�Xԯ�X��o=�e�#����P�[}��R�D���U�[Zk�0�GA�b�#����A]&}����ۆ6,�Q�{���4��U�G$BU/���ѾI#՛�w���f����a� Ϋ1��\�{$�b����Y�E���܄��p����ê�����܋ &�!�v�?�	�Rs��>|K���zA���;���/�c������e������(��r�1\4�-��.)�{��eo<G���Q��6�d� s�5��_��ܳ�1k.~����)���M�j��)�.4T(�y��" 欳-��g�ʃ2{��%j>�]d	MQY[I���d_�Ӡ��
���.Tg2�� ��*�2�|�Bl/I'8������J��Ձq���t?�ر�����@�9�W ��.뢨#ղm�-|��ZY�58i' E$����Q�r�zB1xW�;
f���!c���.7��kY�1��⟝���$bcM{\_,��㎆t��Q���rpS���g6_�, �bh�]�`����@p6�V�xF"z=��[u�g���bA2�����#P͸�ttX��W<��^��+�qdx��X"���v%�P�����!��KP�i��{�]�U�y��o�-T�ظ��mnW�)���N�k6��oy�����Du�F�5Ԟ�(	���l��N6��Ƣ��8G��<��H�Tۓ�G���ۼ�\x�.6�5��xn�#��4cW����e�3���?�@:��E@�R{;�˘AUC	�� ��>r^#���RÄp�_�3h�W�E�!�eo���e����7�1��|�ɽ%���gA�>Yǈ���1 �9������g���۵*W��L� ����U�F3z��!�p�����V�ڃ��V_A�ݫ�/-\X*?��Tm���4l�ܑך`���G��Z�7%��.(���YN�#�Q �[]�;l�+C��Q/��A2�������DV.�Y_��E9����	�%Q��~��Vt����f��l͢z�o���m�Ák�3I�&ĸ�.}R��\�ڼ�U@��E(�Un��)�W�2_�7�:��\h���,D�pZ��B-	�T+��pRg[�裀I�K�mMMx�f�X�H���,�.4F=����F�(�F�֊HBziU!G�1������Vu����S5զFb��1����/y����A�1���g�:N�0Z���=�9�O�jg�����=P�Uyxv>��l��ޯ�PObޕܤ��͸���R#AR�M� ���D�\	ď��vb��҅����l������R��W��N��&��%����"ؑ�S2)��5���֨'�IPa)j���J�ic� ��'���<.���A\��'%�?�q�YK�;;<tKt�dXY*���"���}��j.z[�i?�hl���4|r�Fz���P��Ohd�֧�]�Ϯ ��i�}1:hNs����C�E֣�(]�D�G������=�w���(wnN�6�Z�֑���.H�7��Dz�
��B� ÅD�=C���gS;%�[�iE5� �O��!�^/�-�?���GZ�^ ������H����n2LG����/X탪�{�»n�q�����H ��;��в*�^��N�XԸGw߷�������zH����A�SaL��>K����d�q��hI�7.��i�їɞf�7�K�J&z�ݭ�J�L)hq��4^FD�����5Ⱦ���YN~���D�\CP6�.�yѿrX�?�?J�� �Q?J��"�2�ߐr�~1��?Y��e����S����F�H�.�ƧBk�+8�bC��fI6� �B�R玍������)�oF����q{P^+�^���'�o;)U<�\^�ƺ󝎤AŎ"^J�����m����ư��v�0�\�BN�6�)�<��m��/��lޤ��C��2�6̞���<��b�i��`@��n�Z������+�=LR�3��g�dY`�#�~���Y�>�������G�� R9�����K�+��i���ퟎ�½gz��e�j)��*�9��p/
ZI��g�M�y[��X�3�E�b������ 8�/=�cdA29h�V���x�M��G�
H0s�A���y_o҆Xz��,����&.8����&���=��D��}��o�佹��Ѫ�|���%D�ܟ�I׮���㬣zȦ�!����at�w��N%�{O���n"�%n8��C���b���p�]�5�R�v
�Dk%���60Ry�)2	����C"Yl���^��}��B2���҂	}%�>nr@��?�-4Q�<��zt�V1���6��(_��h0��8�׽)��� a�1���,&��?���4�00�Aca�a���fN�/eo���z\e`�2bO%w�pn\ i�8�43['H�xZa��u �0�( �}�����J�;�,1hu~���+1
M>1�.Y�.%g�U�� �'����R�e r��mԇt�a_�8[��ǸU�o���>�1�ˠiRM$��
x�՚�|��OԪ�[��uhY���A|�(����MeY�%M4���vd�+ ��%�@/�6�ofv�fGL�+B�?�CW���a�q��y� ��M0�F��p�M?s��܀\������[�Ϸ���L�֢t+9Jp���+��?������&��sGV�7*�<m�n��-bF��QR9�2C%)a��S{����y��~�T3j~2�qT�I��o
�r8���$�o�m���C7� �SF��{�M��凁ި�Ի��V	=
3O��3���ߵGgO�t{��yM��?�QoED_����.�V�������5ӈ�r���O·���O݅?gpt*�t%���`~�EY0~p��^OݞsCm��'I��@2�{��J���H錟�;t�P�P� /C�]Y�� "QG�������On��T�	'�=7���V�����ǅ�ך��c�]u��M�±���K'Q��z�����O_E2�!O�8���%*ի��e[��m�b�$�}��J@xP��|Fh�i� �!I5�tW�d��N�\*�v����lLc�V��[���%e���'�9��m�?������mNN`Y`�ϡ�	�,m��mXW�\{�XC��'��?˙L͜��w�?<�&0L3@�y�}�#M4}�E�j�����^0vP�)�&@'�*�J�!.�szmke��~��Z=�&K��j���g��h`��g����}�i��s��t��<�Y�&1`����U�F��5��&0�{:�(�^�h)$�o����i���\������N��o�	��K���;TK�ro�6r{1�W<������Z���PZ����~��k���N|,��H:3��X%} <��m��> �����dT����D3�,�;�?�; ��	����J��`�*u&�0���?��H����g�B�~�ܷ��s����l�"�����y�<����f	,����e�'kֳL���T�#���s�c�X�Q���C��ƍ٘�߂f,���c�B��)�F��_�ߦҘ��b�j�����5Hh. �v��d!0�
��B8e�9�������f.wa��E�������@��[8
9
�U�CS=1r���m ��UF!�Nl׀�H�D;�9�D��Pۯ	̆ܦں��.�.R	��w!�+��W��ߟ���w/ے�,��a�M�S>Ѐ�z�K�w�;K����:-n;h$��r����&"�I��@Sގ��A�!�3����?q5��T�{LX��s�7����w#��)>�RZ�V2z;#�l0;�l�T����p)�/ļ�ɥ�� �#�	��L�y��rlB�ŜK�˫�e���)�a��^S����,B�43;�v���^4��G��"ВEZÒ�E\ �'b�Gƾ�
Fw�Ljؿ���Z�_�?>ٛLR1?@1��N�`�Kj\<������]�����U��V����?~2��7�*a��5(���}����`���G��hf�ǖ��gD��Vq��lN+����"�	n��V��'#�m��^vD�����n�����V�mD'1엑�O�>D^�m�����54.��D���ۊ� f;[���HW��c���o���ܴ(Nr�@lؤY:�Pw �u'�=���� F�@Ѵ�Ƴ��C+��b3i�<����c_�X���*Ej�4O�c��|�O�����m�cˬ���٪A4�3����Z��H���2�~�x̽^��W���Tj�\ct5�����_�c��_�dF� �[��waIi(r��M���0/��Yä�XLa�TY݅R���mڇx`;$*M���e�1��4	�^j�	.2��I���9���netC�$� �U�2Pr�FO��������`�)5�>k�T����Y��Ʌ%��Է3��iB��ZYB�oZ�5���nĽ�8PbF����.�ZvU��N;}��0#��MV�|-�h�;���Q/;EOK
�$�V*��inDt g����9�2~?��B�I*����q ����$���&�27�L��$�I�-�H�^�F-���١b0cƣ"{�C�~�VsR�������
�
W��Օ9��wf���־.����ό=h�<��ġN��S�����g�fz�R��bOCF*��֔�b㚺����A�8ć��4m':��3_�]�`��x�M�[������ ������$2��A[ϭZB+oghq�S���������Tf�k`�mc��u�>o���jܭ�K��Bw��g.�)�4���R-��?6v$����M�/�5���K�ĉ��z�̚���ڮ(��u����#^�b���i���߈*��|8�;Xר�XB���<|�Q�߰!�	Y�8�լ967wK[[ #䵿�Su;_{�>~7��k�l�4/�6��߆��#<3h�|��%̪,g��'�n�UVJnmǎE������A��	������"7kK�)?��d��s�]��2tǟ��=GQk���0|��/d�gL��D��xE�2K���3]&�I��$֋A�]�܎{������=��V�h<YH���!D#�H�#��sQ��i`z�fB6Y�q�~񒠄�#Oo��g�?�8��[{�ܼ
�[4S�!$���6�W�b���\�}��bgjAtd��#�|�_<1p�T�e[%���i�B�V�f\��˼����45���J�{W�}>�|H�<x�)��M����	��HRP!��{=�Ē�Ж���9��xW��CBͶ\�҂�u���)�1�8ø4��c ��c�NnKAF��wo�@?��K���̠[Ĝ�2asI-˴9�&�l6~�
�O�>i$�DU�g�g�<	f�5~����� _Co���V�i7�s��� cd��������z���Fۅ)���۹R��^�}=gj ��!Aږ��$�^���A�	�4v��!����� /���C|��v��>6Έ�#k�f#����Y�s1\����FUx>!��j�#�53�1��	<�>n��w�f�2�>CUFrI�E-d��	r =�5q�1A���˘����9���П	�/�� �!�T�O��J5q�հ=���
�L	}��,I{�|���&���4�՘��a�K+�������K ��s-/��@t�춯&H}�\�'����^(u�`̤�Rf��������_�^w7�tȨ�e����ڰ���/�������M��8�ÿ���M�1ƞ��c��:V~�w��!)Jp:��֍ڌ8�Uu� �!�k��PY`�49����,b��2�w���Y�i���	����1!��Q��P��^B��z>��ےWi	R�!p�R+G��E�*4x��I2�Q^��6?��'��5���;�R�DS�����o��.�"�l*<�P6��ϝm�=H�D�|�Y��i]�^AzV��TC�fi�7�|e�;�-Z<S���o�i
m�$�l��AP�nx1)��Q��m5,8�!;�;�y~I�%N�5��:�����雗s������>��axpO+��k�`H���$�I��D�uo٘ߜ�s+��J��_��-��}����ԥ�����]�	�$h\x�ͥ���
�t�XWԅ�N�&�NXo=!���������8"1>z8}�~F�n�9e�Q2[!w��[�����l|�bN��e#�ǇS8v�������hm�q�ٚuG���cbK�om��9l�VC���´li�*���)I������ڿT���|h��G��S�eϣV�|�%c5i��Me~��y���(���O`FК��f��l���à'�͜���uV}��,k��������3�����a��^6j q��Y��QЙ�K1���9���9{�G��Da�=�Ҥ���.y��:K��?lL\5�t6���~tE�����8����W��+�3��v��l0>�Y�%��SNsz��!���Ը���,�J���	�b^�@��3�����E�U���]�?��V�����8A$�SE��c$F��N�lp�Fv�� H��Y���Ӟ%K{|7#��iq��#��Z�5�V�'�m';�o�����zRr׵��?w
����7�_������t��jߪ�=Z	�H42?��;���j���\t�]�קy��G���/KGs�II���<n}�0�
W��_I�)I���iq�(��ڋ�>��T��� "�y>���м�cڊv/�M�3q3~@N߼J��v�\W'� ��,UU/k2�r�C�m|�FWd�p��"�`�EB�A\�c�(�ym�:ϭȵ�~��N5�d �"+j6ؓ�C��n��s<ZG�������b��	���k�$Z�I�|
�m�D��b\ �FsIq�t�}���M�߉��i�<��W�61:��:��E��z�CV�_�#�Y�@�`��Iu�~��VH&��M</d���"�yk�>_�<�`t~F�Ң^��$��ĝ�WR����m|W��� �`�fڄM�s�t�*VON���ľwuq���f��TZ�����`�<JitN��<J����
j�tF7pU��WK?ҕ���.��� ����끰��d������?hDFaŹ�㭖]9���g=0��C3��`���̫00��Jo}�2w�X���O��5.���&�Zr��@����{w�Āp%�����e�H���Ε�3�/��e㚏V��x����_,��5N'�[��eE�]���unV6�gv	.��d	�Z�����7�Q�%�S�厱���-�W��=�������?��O�z�����e����`%�ؠGɏ��������r8j��Q��M4���0����=ϩA���{vE*��5�dpY�m�`��~�C��CMH����2�R��Z@!�׭�B~=�1��h��,ܩ���y�: �;�ɭ�Ώ��7�D܇��&���lw�����7��c6A�6<���*�h�NY�*߄
R8mMrB'�`4�����1�K���GZcSׁ�_��g�pPS��##O��*O���b�c�?�F&���j�������GoX#� ��`�K�oL�=�hSW��	ӟ�\��Hg����!�P�<m�JUUL2ҡ�0~��ũ��1���
Lp,u+ga�a�dь�HJ�;�ձ/��+����\S�+i`'Į����}��
�e��D� 着t"�+'��IF9=��i�F�^T������Ε+<M�_�Rw4k�V�Hۮ͚��1W��9ݜ*b����*+0nt�D��+��+�U��,�Ys!��:��Gg4�@��}N{�H!TC~�I���x���t��m]���ܶ_�����6(� v����a	�i�R�A T�ӓq8,NS<=P���gĔX&��8N��}���ضa�կ�`�a��(:N�����́��A�B�՘�}�����k�S�.+� �,��z�Y�b�"gd}��	����m�S�T9m=>����K�]�Jg;Y�|�k�K��h������n���x�_|�ӂ#�
ًV�^�ޗ�Y5�N)�	
5���ىS���.$ˠ���4�a�:X�Eq�`�����ǂ��)t�q����`<l_A���,+?M,s�ߴ�_�@jp	w��W� G߀��[<������kb���C���C�fQ�G,n�/����W|��vn+a����n�j�T���Ć���g>M�@�+�+[V�@��8Q�D���W�p W$������c��ܪTS�T�eyA�hr�T|]
�CD5�o�lS���ݰt�koRt��{�+L���tkN9i�qt}ok5܎�K2�b����~�S�}��q��g��>y([��;�e'�R������j�a
n�9�Q>�b��O�Fv�~-%��]�UD��J��6;���'�K0j E����@���=����s���j(�$5�b�Q�t�5i?�2%rE&I;���KՅ�7������}N�P�o���wtJ�!u�%���&��v�G�\D�mH[����dJO��t�t��1������k�@F\�������?�o��L�b���_ʄ�ю9|A.�b����xV�c00"���p��%��.^;�#�oR�pX���tA�J�_&��*���q���H�3�x>63�X����5MB}獬��P��p^�>$i)oD�]��ZJ�M�1���fM���ku~E'��f$S����q�����oӪv^�u��ĭ�}���Bi�e:'�
e啄����,G_�Sx�T��9�Ed�Ku��CI�&V�0i�n������)��W;}0^˟���O�4e���\��>���{��5�-���6���<�-��^:�Hޒ5�� ��U���Q,�7�kC�d�'Y䧑G^.�!��xʞ/vI��fR���4#�]��z��������e\@�eμ��ǭ��)p��/Y<��Wr\�!ɛ��JQ�tF2 ���Ū��.Z$����֯�ܢV�-\.��wJUYm���v�b@��i���Y:���J�ͯ�X�uW���i���[��������qd!~*�~k��F��Ԙ<9(��t�{�$�½�����n�30��8��{��=��3���/�Hg1�|A�b-�B�(�A�zu��^��z��@�W�r)����$c�Da�;����v�aE�_�y�{�.bE�2�@���I%⦞���3�rU�&���~��>Pa�x�� uEW�2��%	q	�v?�.��Ũu <�ey��U�k ���@Ƭ�-x�R4��̨��M�3�b��c��h9����R�۬��H�Lr.�!�x��C�'��e&=�N�==7�i)M@ץ\������<H�xDdR�`�Qy��_��KӘs7�a!|B*D�</!Jw�6�:e��Q���{��6.o!<9��}�wGf��pI ���t�w��A-e?��O�i�S@�S�2�U����;,�:��yz��'�}n  $E��n�)�N��P����H?-T���<���q�A��w6���S���E�
D��3�N�����u7q��CQ.Al����W[�Gpct�/Q�H�����(��� �/bs]v��z&/�i�K�w������u���'��H`�N�Jd$F�+�@ō�@�$�K��߸�bK�F~D����?��XВ��� ;�Kٞ���7#c�iʮ7�1�R��0K��Q��(7h��[h�%g��ی�SQqk�+L�����?�
�ۼ !w1���
��w拦�ǜ�ͫ�b�"'uL���z�!X��vd��0�xD7�Q̱��q�?��l[m���}�^�\OY�ײ��l[Ls�vE%\2$���T��HV��f��[���BOxj�D<�<��2�>�[qHPz:�B�:���
�V	7>��͍..ֈ��gg���t)o����*g�ڴ�}��B�:���H�:��U���e)h}���������;�,�rf���0��7Z%���&)���?���_�7���v�fD qz�3�G��G[S�Z��}�����B�X�$]�ݚ�Ѻ�4D)h�w�T�x1L=	�,�=�Q��*�@ۄ�UQ+��B��ܻ�|ܯ�ȡ�` �W�e�@X��U@!��X��v�������%{�;:pOŉۋ3hG��򊒔���MM�)f�u�h���O�*{S�����֐N{�nۅb�έ���1f��b�Ʈ��:f
�?dֵ�8�@�B���}��3���I�kf*�1q(I����v5
qO�O��A�\�!� ��|X�?��?�]�nJ�w���G7J�4]SP����u���,�O^�Y+G<��UZC\j�.���^�����`����#gy�A4�F�by��>g�\�LO�K����.WG�k�d�L�Z&|!�]�Kw�D]�����3x ����蕾!����L׫�~@�� �h����w����O�P��W��`ȯE�?��t;���Ļ q�#�Nu�a-ct�n	�}I৊	��H䎹�S�t�����h����y�%
�3���%�GSш�K���}M�k4��J�,B��8w}�0X��/p����pWp���%��3:� �%�W�����L=N:C�d�����#��g4)U`^�+30g���s'GՃT���@S�b���_�-㭐��m�!*w��7�X-Y��d	&�9*΁5lL��5�'H���{����U��}"4ʿ�Tw1��%�097���&�� �C��`�@���އVix���V��B ��m�l�����i��v�1��L�7X48�z���u2u��E�#���r��k���{����a�8��c12�=/�ˈp��6I��Z��h�cf��+:��z����8�W�Vq�/���W,�����
ۥM�$1���~�����p� aJl�2��bo�>8��
��NP�rP�1���i}��^wH%��Fo��9�jmT������T0�!�~��J�Zv���b�W]��-���b�T��(��0(�5�D�G�����&��9,+>W�' � �n��?N�e���A&��-#��|��U	1��J�\��*?� �U�X�����R�1��mL��Pem3?��;��͡r��L��FQ��3n�Kz�p��浫�i���J�1���h��n��G[4M���d�B�Wb��ۧ��P&Y
IԨ#
�{8���)��-�G5�4���?yc^-��t񂀤;Q��E�}j�~�W�I�P]O45��#���?�y,��|Q�6+�6��1�/T���f�	�����K����Ž��\�e����hx�f��h�1��
�2���C���ϗ��{I��镁 ~�gI0:��I*��JC�92��~m'3,ۉ�ߏZŀ�V�}�x�
�����yNs	�Q���F�GS��M�J���EݛΧ�����e>�	���H�I�4A��]
w ��	�e�b���H��:����p粴v�����U���5	��M���.�<�Ya�Ʀ��jb��>qo���+D{vgۼУ���6\�v:e��\�ޖ8�z�(<x�����JR���H��0^5���ʸMNaoC+\��2�j$+K��I�n\�{���s�m���_�"�NI�j������!�W�&FHn�q3:m�k��|N?{�D��3u���+E�y��R�qj���_U������=��-{U�#�l��V�{�M�cd�W�� Hj�&�{��.�5�)_:E�8��k���.�8�a�a��TQ�n�����`9A�S�m�xX��fdaPn���g��k�b�?`�>'���E͉x���IV��w�"�Q�YZ	�� $���`f����on?{�fK�����J(��j<��K,�1K��!�8z�;%9v�����<3�v��j� �q�wI]қ�~h����E�=�G3�u��~��(:H:�n����(�IҍeUh��Ol��hp^RKl�!r�ZmܺHp��A8��F�B�ǾbuE��@���f"����~,�m��#�7�.4��n�|��]�-�(�+s6d>"'S�/�e��q�O��*H"��mD��o�v����zչ����s����JA�*7 ��/�nJ\]�Px��d���dm��JQu�yQ�p%���o%Ͳ\U�^AaEu �<g�+�нO;�u�1\�^�~@D��%�&DL�oi�8\��ל(�[k ػ1���FG)�XQ�ǔ�c���:5%
!���F?��&�x��sK���I�G-��zS�~/}�@���7,c�.�L�{,n�$�A�ܤv|F���h��:���mi��0�le�~1����6e��N�_��3���D뇠�"pF�X0*
a�`�hq�]ϛ9������D��0���'w=!�`*�eu��aթ���f�����,�4K�����j��۲��&�l����Ha�e���ʻ� ��H�1��òU�-&�����r±Гz�ibb�2�8(r
��;�^�q��y�Xjz�z!�d�/�1ȞUW����D�`�Y��� �����&�lu-����_�*��ü�p�V�����O�ǭ����>���y�t|���q���h�j]C��n4&r����h���pO���c;ۚ��HZ���2٢�����Hn�Bh'k�(T����N�d�8�d��y�N��%�&ـ���z������tv��1�|V*�m44���%(l�	�o7��rt��5��V�^|�b��E"
��$��H���qL|�P+��9Q5",���AΆc9Ŷ�רo=D��F"��9,�:�* h}4�(�f�W]�r��NW����b�:%�F�ᓣ��k��X-l������
z��u��
��P��L����BK�F!�,ʚ��ʓ�{��O-'%��:S�+��ذ���BI:�۴D���v7���il&�莀�ʳ�����o�]�[�D�ݟQ�o[�u�8|>EР�Wi`~���_]r�(f�^��6֮/���I�����
Ӣ#.?����ѹ�jF;]����$2��@3p���V�!�0���?���������8�L��6��ɖ�pE�ґ�u�v'�
(��8��Fn�8;q��o���
5��ƿ[���I"���0�d��bc�P���J6ɦ��h
���k҅��DY(
��SMyT']�I����D��}+���z  ��ʺ��vy%�	R%ʯ!��<L��P�� b�9��I�������a٦���z�G"Ph��آگ
|5�kA\6�g!�C}{���N�&��m�*3�-'VR���
�;1�Y���o�'_��b��~�OT�󆒷c� ����p��N���4�M2qQ�xb"�\)��e��o���PȞ��2~c5p �#��=%I���=�1}�|��[�:~�և�o�z���Q�f	`̤�÷��Bc�Y�4u]�����%����d�GG*v���1�1͊~(�Cq�F~0�(G�'.� ̋���斨c�%����|�Q��`�5���&����l��q��� ���<�˕U'��i�U�uKc15#�>PR|-ξ�yH_=�U�2`�f�A��F��M��D��2��|��t���DHY!Qj�$c�=pv������7���;�v�_h�l�N�cUUҋ��;��OgЧK��쥓��K����)_�����W2���!v�Ba���/�2�8q �$~���ޮ˗���z��≮%�`�=@+X.=ߵ�w��]�T+�����b�v|88;�B���4��N����+4N����Uü6�@�k��;�| q�K��_eL3GL�p̑��ڞ+B� �R��X���/�U�`�|�~�I!n�63�3E[��onrU�9�&t=1|���@WZ����}�P��g��T��*�eyP�Gp���ӣ�P��-�n��̶�SQC�ˊ�l����~��Ab׿�0�4�Wӷ~ +^��n�0�yQ��s���F)i�ח���<$l��HtX3��6d��C㎵LX���JuE;I+oEaغEuH��Փu������ԛDf�cLh�Gp��l�q����8Y�{	����Sa�Mαs��P�'��D���s1H1�O�b�H��U�����<��Q��ǳ�iY���e�-%���6�Nl1�#�2epx��8��'SRtcr�-?.�,0֝�����I����w-�C��D��0��Uԯ�n���cC '|p�Q}S���k��uƩ�|���X#�9��3Tޘ�F\TS��sH��u���ٮ��E�Z�.<��(�!8s?\�D�0$.���� 1�ys6��Sz|"�R'�Gn�Wd�]�~�:������T������j-�F��2,����r����P�*��\D��M�U�`S%��������}@������ؓ�ڊ�'W�O��9�����Y�'I"�q�2l��q9SN,�����dC��E�xX䲸p�"u�u�)����T�@���Ց���� �����F�[��Ek'xs2����0�&*\��t�K�R1��.�K���̿�uM���o�yV��!�y���Up��iP�Kz(��G�tE�ov� �:Ëd�%�}��wA���]ݲS��ϻ���a�[��ì�?��"�"`����^D`TK)�n�M��"U�Qi>���X�HY	T�]�%P�7���3?ݔyh�'�<��p�\�bj�F�e �����$Y[L�Lo�E��#��C ׈��I��N��#�k���t[��@Ʋ
�������#�b��k�3#C�/��|�`Of���Y涄pxB9�8PU ��4�f��̠T�����L�+�f{�Z'�%qej�򃴷Ob�.��H(��Xc�&R;�C@1�׉�NB�s��	�IZ:&x�N2`�V��)�D��}�Rz¹T�� 0�}��i�&v\���#0�k1xS���C29��y2�H�!�}������� ��/��VL��ː��r�ϭ�E!(~�Ͱf�i?sGB�{Ϩq��a}��%�|�"Nq�����J��g*7���r�I�e8v���"w#�RLHU2��١P��!���Q&���L��4NQĠ�ޞ�2c�+�R�TK�9Xm9·�~FZ�K? ������2�|tIe1��!{�SC�'��,��Bblb�aV�B�.YF��y�=f]QE�5e�,�9J�V�O�����G��wcvC�hV�%���_���b��9�W�e�
�mx�/uch����D\)���c��	wˊ�i8�E�	E#���ŬI>�R�y��rh�[�&)7��u�vD��	�F����($:��kI}`�n�]�_	Ӳ�V��(D�Q��꣒��f�˰����	��TڊβHF[�%#��g��d:�\EEN�M�x��0�]dbɭ�|i�[�1=&!8D�?�S����^�}�&����ŗZ�B��c��:$���4�,7+B�/�ȆX�_�e��RZ$�7���(�vQ&���ӥ`Kh;m����j�)�B�4Õ�o�ğ�ζ�]�c���
�LI��4Yĕ�*6f3Iǟ]���Zqq*�-ᇦQ����}ֈĂ��C����Q��H�ё[	�nc�s�(�+Z̎���+�a��By�#5:U-;��M����mc
)�.P���[%)���k72�6�JU9p�_�!#���4d����`�"}"[)���4��ԟ��6����������k�	����vA>��rq���+
׈�8I������n�u�����A�$�@���!����?]��v���xj��T[?P���*���R��$�7�IC\�8�h��V�r��[$��>�O'�[�.o�~��)\H�e��P�����:����cޕ���@o��lwv�}3�6�K
u=��G���ϐ������ R
�.��Um*��%��rB�#��ե^���R3sۭ�į�	� ��9�G���?:��rK`��@�ЄEzZ�-k����
�L�]�)�������[e��8SPĩ��j�k*�;N�r��Z�C"����[�uc;F j���3wD,]rk~a1�!�2��k�r�0	����D��~ {k2oҔ�nuX�5� ���Sb�lО����z����emŐ�v�E�Rv�n-�d�Jf�E��G7�]�.��,z4���L�n��^Qt���fѦ��5-	%7��QK�]Z�+�P�x��l�t���{�cM��P̿��"o��'�Z���4^m
H�E� �XX�� Ǉ��o�{�Q��[?�e��4�=�E-��1=@�م�L��[������rE���3ѣ5����e5
��c�!|Wr?��6�#<�׾a�ޑ�]�:�8�?�U}�e1p���捛�����&Иg���ء��8b37��� ǈ��2T���z��9�]��J"$ܑ����.�'�׫�a����WUcǨ�~�-��n �ɓ8l���; 9�¬�0Hg�/��O�o��έA�����)�Vg��恵,^���-�qy-����3�)���cLM��Y*�J���8�Nz��t��*됞��D,��ޙ��~�u�2}F~ݺ+�p���0/�_�?���)��;���tn�|�A͕6E�U`�A��|R$�M�TU��5��wvh��=[�0���Mk;ş���r=��P�<L�c���ϯ��_rں�\��q��NK�xo^44��=7q�/���8�Rjz�Y8��~W,�2�}�E�x���Q����{����/f��az�O#V��A�"��$L:��N{�k�ˆ��Zx�u;|f����8�%ܿ�d�R�._:�����!C�F���U�E���/`�ް�bn)#���mj҂7���˭���_�.���{v�z>1�h��Y�� �B���׶�&lY�}$L�fx���K\�埗&�1]�ޟ�u/lz�B�&�l���cǢ3���T��4iJ�bz�8$��u=�3'�����☝p�I��7����!�&z���miү�_�"?5F����������FE����2}�Tc��'���
��@u�I�4�x�^�HؿDY��Ţ]�m�nM\B!�������
�!v�w��,�s;D���?�5�U���Z��Om�_� 0{O�k��8�"�Bz-��?���������DR��Dk�t't։�U���4؝.�`jX��Fy,>�|�4�;s�]z�����	�pќug�j~�߯�S"��/�l�����킏�ɂ��g+ʙ#�Zo��m/��Zz@ڐ]����4-���9
-���J���6��AUf"l���ٍ�k�j�H�7P��8�<�R&yX�ς���$������Xe �����|�n�����YF�$�ֳ� s-(��9<@!��q�٦��g8XG;�~j	`�fXHf��*����W����,x�A8#��#��3z��R�[���� 	�$�W�t#�?��5ӭ�O3�f�5�O��o�V{�1e|�"��wy�GN��13�1���s��
.)��;�`�*�3�M��!�5���9���#�����ϣ�Ho�*9O*���X5��F��D�yѤ]D��G�����'�{�A��v���p� ��PŸ� �����y��IA��ϙ/���6vHӱ�D�������̓i=%gPZ$C@3)�Ѳa����P�%hh�k��K2�:m^���EtS�Rbk��EK�e�D.y�jfE6�)���'K��w��|]�vd�&iT����9gW��>8��g2��T�fe)L��)&ވ���y^��9�K�Ќ�Ҥ^����eMm8|q�$l
�@$dt���/�ʻlְ���1c}&��9Z��Q%k?+��er��$(�#�*ݟ\-s+���Jë�WFS�_�	��W���R�P?����cv���uم߈u^,�ݾ�>��Y>���s�r��,ɂSy��zHқ����|���{u⎚uY4��ƺ���.�Q�YA�dI)2���_8L���	���CE� ���%d�2�P7��bs�\4;�i@��\�cg���Ģ�}��Mqpn���c%O�#�����ik�YP���zCR�I_�.GC�+�]�����z�m~�E��߲+�N�p��j�+�#��	�i��0ֽ��!��YGĕ�O3�~���y��a�/\��^m�
�9�)$2&�NY�}�%��3�hQ�u�j7MV����v����E�`y��`'��0�V�P�o؊�#b��S��F�D�+6�?�X>}��6�����q%�U#|
ڒ�*�ѝ�A��Y��9��;?g�$M��8V@��@杨0$�G{�f`���xz!��2u�n�����^�����ډ����%ۛGBD�S�l��0�����Ι]�"��n2���Rر?O9���r���D	��mq��k�)�~��4Y�U�bbP�,G��ٖ�@s�rK�]�K5q-ɲz�n�b�{��4� `qN �hh�[�
�O�( �6�D7z����Y@{U2nCm���1�;*�����7�f7�>
b�yP��Nv�����,�k�ƙ�:�;�ͮmF]m����X: �X����O^r�)*���kO��λ\�ܰ0C�"��F�x#bP�Xh8�ŢR89$�����&���3��=sUtZI�bl�����D_�>7�n�����!�� ��c��z7Vo>#���n ��������5��C5���D�R2ĺ�}�'-Y�~%����H?��� ���_L)?v�c:^�M�D�� �Ϗs���ֲ؃b���&i/z�S�sϾ�[��?g��F�:��$���V�=��T���X>3�˸�G� sg�:.d��za�wӨ7�tM��K^�)W�!M)C�$oh�9���J�o�j����g�B�Ә-�1s�"'�(S�z�������N;�#������F`HR�+9WfE񂴠 ����ӣ��\��o�DpJ�Dt���#�O�M(`��\�g	��N*AU�Ե�&���3\�c��S�8��^1�y5�	  h���z�-��n?3D��<4�l��#^���Y3O��XL J_�m�}N鬞�{"=b�â������T�G@X_�|E��ԝ`�XB)�O���!i��Skj��+��Y�֖T9�m3���2�r�-�ګ(r�ܲ.��s�;�o���+{����(���/{RN�b����~�T'��a��=���u��ѵ����f�&���r�q<6°�n$L���,!s��L?Q�9�Xw�R0�C2kڸ77���)���k��%���� ���&N)t��� �����J�'J4�%�&$�_�[	���,���Ή��+�)u������0y�������l��w~�����+Q{���2��
&G�5MZχ�7v��Oo�M"�3n�U@:?{����$��o���>���=��,}�7P��&�{
[V.B1p�w���SK�as��Jbg_V��%0v�s}�b�XY}k}�K|L��G1P��v��
���=�E	���}-U���$�e2�q�b=��sy��ړ��l��I�B�v_@)��P+E�z"8�'l�F>�?��Av��da>��E^��	H��������Z��Z+[5)0�̆�Po���|b� -YN�?�7��8�?͗!齁��U'1�C��
%��q��߀��ֲ�Kt�
�+`���m��;���؜�ן����P8ʏ<-��+-oj�� ���3��~�I�uv0�\�4�B��9x�ݹ�\^R�&q(@��g-A�=�8���-��h���=>6ۢ�&ff83���+���h��,��p?��漏8yn&�G�x�Н��WIm~��m���ca�%�3P/8���
X}��s �W��)<�>��(j~���a�H�n��9�:��2u�$�'�C�*��H|"/�ǯ�=J?!��� ̀f�.�E�
=5�`��m	�&@�툊r/�����5��e(&�?)Y��|0�Ea�����P��&�B�L��f�
aؑ<��M�$�N��zڨ���-37�|�*+U�B�al���L7+���g�6����OS�}�vk�ڲjR��CAze���Lǻ�0G�U0�bR��|9��'+�r�#��?�Lp�?4n)u�s�vbɱ��=N�6t�@�n)����.̾��~CM�]_L��oJ�c���t'�Ҙ���o��\�NՑ3�\�礞[�1����8U8� �.�1o0ěN�E�z%�)"$�7y��qW!ܮ�1\��yD'�����غCJ3���Ӟ���1��6Y)�a���j��N���C�`~�DQ0�0�YFB_@<p�x*��kY	���\1����T�x.j��&�g`��҄QLW���,8I��vuqp2��Y���C+�V=��q����j�!��yD����!k{��0�ܕ����$��/�b�`Z���\P�^���l,PA�gvG��è�4��=w_ܷW��kP�M�������,Eo�z���ΈRЛ�^V�bvGlx�@O�Nܸ�t/%�]8�n�#�qg�BA.
�g�W�öN�1,zp3$j{���zuڈ��|�3�����lL�O)���Н:l~�=T�E�h��<�2Bjt\qҬ���;f�y~v�r��7��a�*-�(1�cJ�IdM�DU�p.&�~7C��[�3�L݋R�Cl��1���5*!��z�D�@�����Ak�]=���C9�n(ڎp�Gy�:�Z� ��BCI�gaȆQ�I���4����w}l���2N61}�)}���?[2�֎���]�;#'c:1���tQ����}�C�p7������ ��a�!ty�����V9��2e�QPMT�k`p��Q��B"��$6�����ȟt��h���Zr�O�b����x���?C~*8���B�6��#_���}$\�h-{��M���l\��5���8���*�}y��gt��6�Htv�P{��]]4	tI�����Y���
������!�*��A��|��y9�t�M��6TH�!x�Sۜ{�J����A�Fcgyދ�>9��Q�i�����TC>��1T��T�M��,_��i`,��]��*A����>�MV�Ɂ T�O�>�C�a2u�ؖF�l��O��ThB1>��o�S�����p�q�Q!2�ڮf�c����iuq��h�	�9ݫ��߯���O%sd}�mx3 ̾,�l7�����Ƥ��4['m�m%'�x�s���},/�fK�����#��o;3�$�[ruՎ�����9��I1��G���gǓ�O��-��QUB�N�E},�p}���L[� \t.�F&P���biǮ9��)�i�O���Hc�R@�ļ3�0`[�H<[5s�tk#�cw�)U
̓�;H�Q�G����崎��1;0s��CV��|?����`,#5���L��R��eC�>;%#7��G���e� +B�O�d��ٜJ�_�u�{����p{�_�\N̋�ᖓy�y��	��������72NZ�1M <k?����맘���N���H�W܍���m�����c��V�mj�܆n��\�WhV�ơu�FaqB͖	ů�I<�W�Ή�K���i7[d�淭^<��p#+H�xP�3��\�˨�l��E�֥�Ai���8ι�;�oK�,|Z�-'�17� p���q.D�74G\�P�r9�{�u����#T+_���bp\���&k�t��~�!.FRԇL����9T\�OH\Yf^���@G����v��6��;C��Kqe��v�JY���=n$d��Ɉ%7xk�h�P�%o�)�o��:��ֻ;n���͑Qt\3��@?��-���s��Bv��!גe˕I�ɂ�ob�{j��>]E��CL�;����&yD�V�U�f�>�w��|
\�,�kg4R�'ȗ	V�/� �1��@�b:*i���uV魹!�N� ՟��^jی�Ux5��'m�H�CT��\E��ek� Ȝ
�^�L��������(8s����b5�T���s��dsCIo��;��)�|��[�1��F���7��A��L�مX>�׆��y�+k"���ۧ���9j==ۗc����2��ʗ�=Ȋ�4VD���F(��F,��WT^�+l�H���Hh#��/ԙӗ�T�aCj5������+	�6s�᝛ET�pD� :��2��a�G�?m�����~,nU(m���=�)U$��ћ9^c���)9�����e\6sR6V~9�%\٫��_�i��ٻ� ��/՗�'I#<ĥ���LM"dwhRo߮��w�\)
5�}�k<JR�E9�<�����i�\��H��a���A�VBͷ*�k��zr��e.Ȍ�Q��Uݗ|T��"�ͧ;D�l�<R��x�j��:�����i*fdk"��|�-�� *Φj5���E/�-@�"�T;�_!�����#H#��NA��Xq���"�}_V����c�@*_�e���	jǀ����~��ט�A�1��R�U���i`|����0o��d�d��+$�O��g�w��&:��]���5��[��GfN3�w��3rn}3��Y�T�V��M�e�r�>�x��q��! ��/�<��"e�!װ���q2�GK��h�A]���z��z	}]ċ��	g2�
)��� &������+F�D�q$	$�l�L��w
��90�g����!�(�+���1�%%l\�
V
�1p��8L!�L���S0�2xY����V�K!��R&�Phi�զ�a��J�����[�\'?k��#/�]|ZTkcpX�Ao�][|I獝A��L�D�>�"F��M�|]��5o2o���|��J�ע��l���T����,'��OY�/�^��pN��v�j��DF$�F4���Y��?�P��"��jVҐ�@���<%c#��J����0ja���Ϩ.����%<#T�_��-������^�xW��k�������M����c�ޚ���=�`��h!y���̗ڥX ,䌀@���khm��M�q�h~�<���]d���.!]����h��:pD��lO�TӊJ����B��
��]D�Zᕏ�d�S�к�Z>O�)��������;y�h��)�F�opf�jfC_t��^,�$G{�3���/3c���"����\G���y�׳�k������K�^��B����"'!�Ho���4��X�4��L?1�6V�����C�kv'�{K�a�-��~���7s�Ưf��v��k���G�6pMY�s#�D�͊[�B�$��o�x8������ht��~i�D ١�^7]8��w�8����ʀ%�m��,G:��e4A�tPy7���B�ь�2�(Y$B��h���݉�+�e� �������Y��[>Z��IBZ(Q,;�j��d%���ٷ�+�!~�P���]sա�<�L�1�����9oRh��G�n��<�b�� f��HU�q"_� _],dQ�@md��U�"��B�����V,_�(�]�F�u���p)�����g�"�6���-�'�;*`s�ms�^i��ʝ0�6����g��K�\�0�E��H1���K'��E5u���l֮���7�.�@��&������`3�*R��*������ �_X��CxA��D��(����,���09`<��N@��b�\��=�߾Ji����:�ܰ͠��9BN�"@�V���G����9�E�'�?a}��!�Pl�)���>z\�%�5*n�U+d�D���F�C����W�8UR�<���2�E�c�:�L�j%F�Si�s� �&���ڋ�(�ӈ���j��Y�lY�������uNB��ϡ^�_}+na��J��+��ѷ�;�!���˓�d�t�}4���]DCo	W<s�e㬽$9�c�ٰ�� IWЇ������\%�E�y����g��q�5�e��Fګ�@�������˘p>&߾~� �=�����<���@�����PuB��*5+ƀ��ӵE���q��fE��,�6M[��}[p��J8d'�c�l���~�i%�Bf���ȗ�8S�(Jn4_�X�K_<0�fY`I$�^���y��xfӗ�R�O0��rs�ѡ���J4eq�-���������)�t\�H��8�J�>�-��[a�c�Y������ʂa�b��.5��>&6����A2���ȦLĪ��Ş�PZC(i���OJ���8�8V妨�|�xbk�5�-�,����Ys�LJ����\���q�Q���t�Ϊ}L��a�5̒��6��DyF�#s�S�\����Ɂ����_K���ֺ`KIc��b>�N�Q�B=ɘ�ƨ�ڵ¼FC?�iE��5�f/c0)%&�;Eֱ�Y�k��F��:�a� ����#����	��;L�ҭp��b�'F}-$�YC[Y��&�C�q��5UHk��ǡ��-�O����LRU���7�h�h���T�>�<��*��Ն%^��<_�M �V*���	�\�L9��L�`\�f����R�Gx9�2`*?�p�`�����N�y��W/��s�0��
���H`PFi�8��RBoNDބ>�=8B�y�Z~�۽'�Q�;�!
����g�$�?`�ˠͻ�=@]����r���9OY��	�F[�ݑjq���֡���*��d��Hb�V���0�t�Da�%P�;Uþ��Sܖ���e
6� ����p$c�ltj���D|�M�d���n��eX��k=��qs�Cj�du��!	���0�i������:���m�r�������|�u��5ܤ RY��70]�����uJY'!�UX?����hʰ������E ���XiU*��k�_�f����Lb$0���IjdEԍ��*۷di���b~�;E��Ĳ�j��g�'���_�N��N�s�ܜ(�
����q��w����n&�2�+���AQYQ��0H��Y��>�_G!1�^�lc#��Ŕ�.�j;����{�כ'�j�"4D�Xί(�/��7�ޥ����v|Tfm������	j����Z�$m��(/�'}/�n�O$�?Y��P��Hɯz���N�j��Z,�(���ޑ���Ӹ~�?H�j�jK
h�ƫvp�ϫ�� �8��;i�L�,�ڍ8�^1Ů:ʉ�^G�.h����&���-���ݛ�%a�L���8ձ�d/R�5�J��g*���j��<�>oi�(D9����ޘ>�#���o�Im�1�w�-�
V�5M&O�ThZ��yr���Mָ��L��^��])!�N��D�A�`qm���C���_�b�Ҹl��y��E�gR����T�Δ�s8O�@�K�2G�Fˑ�s��tY���
�����o 8��ia
�x�k���&![룀	g�m�`Z�Nh TPUU	S�g�m��Ic!8���6�R�TCn<� �0�L�P�*�]��X��9c�nr�8>̫���*�\��X2{�{"�Bx��>#h������t��ȳ��p���+��浅�.rN��j^�C�+9RG��-��\{��D�h�>�x����F���>w��)��|=쑞wp��Z���!��U �Fo�9�q��ZK*('��ekz���b�	��`�x���$�]��R1+�r*Бn��d��:>M 1����):����%I������Q�~����,S��Q;hgi�Ƣ$��U�+��O��.���v��/���������`l5�)�����ׂ��c�o�����L�&�杗?`�7lq=naV��#Ξ*��U��n9
�lܑ��L�af�Mp��%���7����E�5:bS�x�,��y���먇ûfH��ﱝۇ���G*��w�1�%�����`->����栵������P����TSѥR�s,df�Q��^Sbi�[7��@5@׃8(��/����Q�qrQvʆ'zC���n�
�9nG��o�� zn%[f��Î$�gY�Rha��\��.Z���Nm� j]���-y�x���Y�)��������	Sҟ�n�ǅ���F�%�ܐ���	�i�~7q�2L���QƇb�yϰ˜���l�O����2��k~��%��)@/������&����m���Hp�=��ْ�����ֻ���;�V�j0ᣙ���7�l>����RKz�`�*�V/G?n�X}l@�L$f���!<L����$A�>	*V9q�X�O�}��P$��$��;��e�
&����y��ݾ��J�ͪ�t.4kLnu�����*�����(���m1��]�m�.�P6@���!=��/u��� ���9ӭ�'j;�c����8�h�o�o%�9K����/�Frvo�o�����j̥_b�i3?�`��9���F�K?PR4t����G�d����
�1��'�z��eO.
��t��)�8�#��*���WÛ�k��2֎L�?3����_�WE?!�&���
٬��9����OL��Oi�W��·7�U�~=Vl}��D�Q	u�g���3��鋾�,��낍m�c�3�Y��N�~�^C߈xx$혮���tE��t�/.Pfv��s��r�E�W/�������b�_/w#n���B[k.���)ֱX����
�;H��9�E?���m��������i��&)����a���F��ugP=��*�#��ŀ+`�D+�r ;ql�`�"]}ٴ�(��
���9�-�"�C�"NB�Ձ/)��1c��b4SfR���.�"h�2e�Z�V�\���kBr� t� �{��/6�FbP}c��}p�ǔ<�w�t+M��7i&�6��,Y(�hO�e�����.^�άI-j[ij��]�<����[1�����f�J8ď�꼂X� �t����vQ��*�L�m6E��	j��R|p�|��1~Et�K���R�F<ީ�|.�0�X�;5l&��Wv#����y�������ř����FG.���3��WP�u6�1����W�=�u�My�
��MSHp'~���6PLRVp]o�t�!yS&,?E��vv�-!����}�,{��l�@J��Ś.�ħg���?"3W=���Ҁ�v�+�]'��s�#{�	Ȧ�.��qK6��/�l�3��j]%�8��~u�7��+�:��)�s,��F^����IF�k���U`8�����bhy����n��$�,�-T"T�<z�l��tcӈ(�\�u�ڝ�n�0)���a��3e�E����n)LV��#�jk��h�}>��YFJH|�KF�[�x`�-QXA� �c�[� �uM�@�E�.�~~�nLx?����FO� H�C'kx�n�F��U,�{�H���H���Hr lzbXGY�9�XC�+��� ��|���_J�\b2�	r�����;x�{$�SQ�֒vO���&^c��Z%Q� ��*�I�[���+�]`3�zET�@(�|��l�ُ(�e�m�(Ǆ�[��3՝XK����ĀKY�f�S�{l]siito9�W�:��CO��4���$�i��:�����4��{M�R�&O�S�u�Dʉ�&Jw�M�Qњ!R���;Z@��>e�ЭcHo��|�(��������ƈ3v����������N����fM���>��6b�S�C'ϾA���a����O�w֩,��dO�>��~Y�٨)m hG��+f!�Sgzre���\5Ɯ]���'	y��: 훴�q�v}x��Y�NG��%X���m��B������4nPM����g���v ��޿�R�X��6k�Nȣ�$� ~�g�{N9��m�L_x��{)'f��M�"���Y�����Z4\6�z����L�ͦn8�C�P��GuF_�p?Ͻ��+=�k����ok5�Y��������+M����*�@��F�(�;6��*�IM%SB�eȕɮdq�&�}���3�M�Nf�/�>_���"97&M%Z9�vyf1�ص�#�e��Y��MW�Zz9�XkT��g������T������wf�/J��f�(�AV�TYI>Fc[�#�]������_��K�D�Z[wP�Ǯ�"mq2wxA��&����x�yS����!���(j�bs����ux�mK�ؤ�Ωf1�($Q|-�������f�!DP���,� <��*+g�x_;�n"�K.��r���z�`�	U��y����`}8��'ɦ�Fu�3B
�K���A�u�Y/��,Mh��0Ȱ۴�}�^�5�0ԕ�|V�䭸�c��H�貾V��������8���J.�����w�ſ� �Pc)�?��> ���|� ��br����%�kP|A�z"��}��Lӊ�����'��/:߉��:��Vc� ����Չ�GK1i�e�Si�&~e��i0j��Yק�_aN�g��Y&�}������EV8���S�a��~��ZB�ހ�/�R�5O& <��:����!��2,��n�vzPr�1Z׍�:T�L��g4������TG���0�����u8Ɖ�bO��w����G�ē��	uCk��*S{�����,ϥNc��:B8�Lh)�ۇ�Z�\�;��ذ�6����F�T�rAS���p�ӊ����+������|V��=lH9�􉩯Ip^Uq�X�n��"�Dtb(
>V��R�/�_ꁐ|�L�';�$�U6�:ɜ��Rڧ1?M��t|��1Q�,.=$wa���|�Q��LWɣG=��`��ǩ�X�{4����i�1����i�/��Y�v_�L���X�������m�FX���=y�h�`�4/���%���C1~`8��H[�W=�M�&�P_������L�^�$�N<\�)`�Fj�z[W�1vJd�0i�Ze�O����8���g��ҟ���Ϛl�{s�O,��7CW������i볎C* ^��>=:<J0�0H�,��Rɹ�. ��ORv��"���n4C���T��vny�P�W��̡�� ��r��Ĭ?�V���3o\x������׻�=�p����դ�/􅶔��w���lR�Y!Nf�U�����r�Y�j��q�vt� w ��r<Ä�N+��}�q��!QK-n,���wu�E�x���}�����(Y�Y
Y8�29��R������9'Y<RZ�y����z!�OW��,A�~�o����"u�I_{Mr j2�8|۝1%vIC�VNE��,.�;-EQ8�إ�.�(WV��"���x����|)n��7���H��g���F����몔qc�ڼk�[�'1�ڄ�b���������8g�ȼ���H���]Zb���}*���A�r��p_�b�mC��ZJG�I��^,^l��a.�IF��If���n�\\����@����Oa�\<��L��,��]��޻�-�$�:���R]�N���=QGL?YzRdjo�eZ]Q�\���1xl�H���G'\���,kdhʺt����������zH���O�F}&�Yd�KN���s�.)��G\-{�v0��>���������E��)��*ܞ�HAj"�����>�nK��@"W$�+���4�`����	b��`~�����ԑ�ZĒ�u���*�X�\/��o�X��5��x��B���E�+��y�#��W���j��#�*�j�z�Y�R�Qjw>=����dθ�P�^��\��'�c����Хe4�F��9�Q�H;|1?�l���86��[�z3��U�V�z�7*��z��P��i�h8��k�S�YP�6��I����U
���b�X˦��A�qR1��ћk;�b����Uvix6t�$v:&U��>�q�7w��.�.� ~\-`a4��;�=B��揶���Bh�A<��� ��Q��D�N�ؾD����1������u��^Տ�ū	�n-(���I�~�~"��,�t2��������f;�E�_̍�"��<O�`�KiL*"������F�?���oMM�fcT
f��_C-2�3�Vvf��@��x���q�Ω�
�����H=���>,f>�l
�ʶ��H��x6C���>���g׊a�p���p�A$r�%�^I�H$~E94�p(=�&������ا�s�B-)ڛ�����4�Fv��i|7�F����V���[��Ғf|�,��b�
�X��ā4�=�g,¦\}�Hc�����n��ϔ��I�54�e�{z�!���S����!�CAߍ�J������\2:��Q�4�}@���{�0dlbg�����Cm���E�4�o�M�~)r��[�SG�{1�|Á�+͂%V�0C�y�E���뺆��rb��w���eG���/�� �z-��]j�e�$?t����Wc�L�ʜg��q�|�\�������>�I�j>�ݛ]�X�AXb0.Ƌ��M����I>�OB��R��m�	�32�g���Ȼ09��Kx7�q�~��_�8DI�RR�;�r\�#Tj�����M���̻Po������4b�8���{�%+��Qp�Q:1�s(���A*F������ѻ�^�����Zq��6v�ٝ�^���TM��#'�{$�Ic�����%�_��r]�5�V��@۪�v�J���u�ed��$;]�� ;k%�v�L�ŧdC�Qӿ����7'��r��Sw�����,J~�Q�'K^ ������q/9���#"��%��)�5@+�2Hl9�8��&4��$��s�1.�d����͑�'.t�~���o�$α���;R��u�t��(�A%����&��H�_W7���9�LTU �Z�E4��J��tK�HT����g�}6K0�	��j��|+��������Ϩ�׹���~ h���(W�@�������s�;��b�8�WIR��O�������0�c�%Ȋ����c��P�Y+a�eT��z��P����� �R7�?RKRN :;�.�*
���Q����L2{-2!��՟��'j�-����(���2��=��>����V��nP�!���#1�0�����6�|U[�t��v����F�@�#���TU��_ۿ�����l�Z�4Z\� Y�c�JzM)��;�Ŝ��cw"2&1�E	��|P�MN�Y����I��3�[����/ ��X�z �.߻�ŷ����SOա�\׶��d��"��:�N�,�\���	�*�k����]�Q"1�2daɢ��Q3姵�j,)9��1�����u&�1
A����Sݮ�������&O���y��� �>�v�暾�v^�}�����nr�R�(���4}q��:P($Ut�Q��)D
Xd���J�S�E�K39�<,R�)�����&� I-rլV���y�s�Kفxe��{ g��+�5,�6ϤU��d^��8:vh�D����$���G���4��/������L��رE^`��(�ƥ��O|�ÆND�_�N�B��5GP�Z������e��T+��ˇ�j(�F�+b	�#b���C0�XT
�1�}�LT��b]Y��5~�&,�߿�T�!i�j�j���!���G��<�9��A!��zr`����w����h<}��I�\Z�X|Y� ��ȡcaŋ��T�k�V����iw�围��U	L���c�|�t4�j�t����,C�r�F^�P~L���Y�'�����;Z�}ƿp��V�0���J%V��x0����_-z���!f,A�_�>("D1�@����/z��"���	=��<�@6st�_�,��P(ǫ������7�+"n#x����Uռ>�:R����B||[*Ţ��".-R�2����9��?ȵչ�8�5�XX��\4Ț�$��ͣ��%��\��3�r�{�/�3x�2%���We�%+�F9e毞sh�<��6�̛ ��R�##J�/��_�J��wg����K="#Ħ�y0	�f07��yا����_:���Ѩ��kף�l�q�Toq�����.�}�������/ʈ�3�]Z�@�5�ȧ_�'��x����^�Am����7�r�4'J�|>���+�ɽ�E�#���9G�F�k3l=�w9=~�]wy�Fa�L�ׂ����ި�#�}�w?��l��!500��h���87_��'��N^�2��klv1T��̨�������J���|	�E~k�����K�����琕�i��6M��Q���M
V�[��q��D8��v��[�^�z���w?���޲�����r��t�1^{'�u{F5���X.��A,1OL]���vJ�Zn㜛�{��_��f
�&��TD�얨(���/�ϖ��#�.���(𯆣��&�E��)z��� ����p��߲���f� �xΏC�d&}+���,ɂ箍�1���[j�";C]l+/6�j��˔�xq�eоF@����}b4ݠU6L�� �#� ׸�1xz�����mm�Y1�O��bd@;��X`��� ݠO\mܑ9X���8t1�+�	[F\��[򏣦�%��bd��׽P��Z�z�H����D(�����µB�M��������0��I%��юT�ն������Ft'`��n�P���2=��=U�n�h��ث峊�<����d�R|�`������U��gϻ� ��8����5aj%�p��R5QP�����:�Ջ�1��������x{ucO�7`=�T_�DQ�7|��ݢ �y���"`U���z�I!{pM�SH�%���p��X��}G�W�FdWhQ��Y+��P|�����gc������n�>Ll�f���_�^)G���A�8�&/U�$G��Q����hkk���x�4�*���bٴv�c�P���p������S�P�ך��?�m�]�����nv)�*u���e��~�c����a��\�� ��5����y�2q4��ϡ)⠙��(I�lv���é�R�}K>��(&�s� �lS`��.�iŌ?
>Z�@�j:UT��=��~坵�J���)ƒ�����m�Rmf��Z����$9.��Fm+�r�b]�In�N>q���!��>^��I*�ܯ=�@��Wm�M�F���n����E	-�t~�saNoL��cZ��篦z� ̲�����h⶗��&�Q�(�����a����,na?*㤸�⦴f$�P���ČS&�3�\'�2pz�ۼ�G\\Ic�G�u��=7$Ef��e69����
:� ����6�մH�h�����/2�,f�bwS�r2q!҉)���Py�.��L:	P/���/ua���|�t�v:����� �����tM�bv+L�0QQB���?$��*"FH:�˼��p������_F�7O,���c�b�����o���?*�wF|��H�Fu�,J��?��:����,��`"���d-_d6�A�W���S#<�l�Z�#��L�"j#l���f�K�'7����BG��)`�D�i���|�`��#]b-�6��~umj.��j����Tp��[��c����P v`������m6�Gh����TdD�+i�[�ڣ�ʪƓ���W�*NDrlvU]rq� KMLѝ�	�6��K�\��[襖���ɸyF�x���+>!���R��Խ�d�$9}���a�=�'*��Ex��hsM��\�궬�3����U�La�8<���?B^�Z���P�&���'�ѧY5���nJ*K1��7��h�4��ڀ$�US���1�ׇJ��B��4�ܼ ���J���;=�yĶ�-�<A�q�tg��ȿ*yx,K��u|6D����`���GM6���Bp��u>�.�F5]^At�3?�PW�O}��jƐr��W7�PZN��� h�c]���t��0h�_�!����W6�&�$�-�s�u���N����;a3�3)��+	��u9�f�̽7�4���ۊg�[��Kt���d򤱷�#��OX�e M��r�@�g��Is
�%���I�����0"�.���GKpQ+4T9�y_��=��%���J8;W��̓)k��Yww~�H�km,1Ԯd|iV�~�<_pj*�!�'�� ֓X�fW��&{����q�L8F5�S�����g+Gk���j�C"��G�V����/�n�Ob��+���f _��`�8��M��Z��+��iB8m��]�8�JO����m$��4�3m��#I:	�ؘ��w�X��8E��೓4����"�L^R���y���)�9�6����[��t��s�KM�"|�A1��`k�<ZM0UjI��q!Z�/ɚ�t5�D���%h����vd���e�x�@Nn͗�Io)=^�P6+XϮU�۱p�˓	%��j��AhG1�?"�P�MG����#�d�>��M�m��L�/�N����ۓ���<���@��AdZm4��P�}>҄.� \�d��W��	Ȋ�AI�P��
��=�
P>
�:\<�֌�<��cV�Ǧ}�R�K��%�4.�\)�FM�����:�]CDT%p��=�M�Z� ��^�YMuVeR�=<�Vj��7�J���a�,|��ɐ_5q���=�%�#1�8X���ikI�p/B�I���;�ze-�<�d��)�&�$�L�M-�Y��I�ޱ�V�y�>=�l��x�KG������,H;k�.E�ܿ��+m���Ȝ�ȏM���vr�U�/�bAc[W��kA�##q��'�����|����Q�����k��E�����p
�4��C���DUd�/t������f2 Qq�9�DۿE�>�*��,�*�sf��5�]Dk���mJ+e��t��4�v������I6�l�d�����B߄�Ȧh��%V�&��f�Y;�%���C�p�G���0
۱�V�ҝcw���tkD�ntbh��+h��qi�؈ �b�&�x8��< H��H9�a�N34l�u�_�k��.���ok���۸-���s≀��e&��f06jҝ{�F�+KDz���ӻ�N%�f1cD6pN��j��;�p�+�&�#���	�qۢ8qX�o>|�_��pu��A�F���YQL�wd+�� 6h�Wr��AJď_�#vE��qV^f�=�r��r��c�9(����?_X��r�G`��Zߴf��t�r�f����n,م�@-�cz$٣4q�[��ha#"<�i�@���0�^���$n<�(��Ј�s�h��͔��$H"b~������Gj��>�g�?W������/�(�?h������=�e$��Ő��O
7��}�{Q�{�1Z�j�tGJ�ߛ�h��P4i	R�����)nwf	�h�|"/�k��
!�mE<+ޚ��I.��Q��"Nm�� ��u�;�9N�I���#H���0[0�X���zMky/O$F��חY�b_�!P>��,Z�<w��=<:��2W���R��P���F�H�)*�	��)�#�E���ߦ�g�LՅ|�������;U���P�{9]��h:}��0VV_��� (+�a��@`�B�s$�����H&ɸ�~S����*��� ��Z�o4srnD�Q��zA�۽�ޖ�ʆ�f����	i:�(���"��VQ�-�W��H{�2w��[�˵y�ѹ�m����LTZ�*�P�T�(;_\��U�cx �<s.0b$�
:�X��y7%1j��%OH��6eW���ϢB�.[�9{�K|Wz�̿S�G�Ҩ,]�)�D	��L�Z-ȴ��6�P��h��P-���ڗ?�����a<3����Zu�wo�턤&j��"I�����*S�{���/w����L���C1D�8jʬh"�8�!����eF��npx3��Jd|6��Pr�������f���N;�$*�2^ڢ߄8�L�f�ޅ#�Z�p��B�+z�2��q��:B/\�u����4A��\L������P�ܟ%߆	���&��Z�(v�ݧa��:X���dMe�����rȔIY��S��&��f[Zl�i����h>!�z�a0^���q�4�Z� Y�ʴC��zT����7���{p ��p�3��{�(bW�b�2}
�8���"�tDKY�bsZ��ԿR�"������yҕ�x�/�L��<�{}\�t^�[�#�Xs~sm�N�i�����C��AH8�.6,u�K�F�ؠz�6H��\���L�*dg���<.D�_WJ��#:T̊nW�Vu�a����H��K;d�A�}����~7笔F��d�
%����w����v�+B(~ b�tמ`��>\�n:�$9����$�.�‵�D�~�u�(�VW h�&�_���R�aOq�UWY"Y%�r��Cn�99$c�q��h�q�dW���8/6���S9�[0Լw�$1���KH�CQag�6�ܳ�7��s,zs��$�NO
�+Hb�(=�D1IA������ak��E�ч�C�BP�퐬�1a�����g�i9B5h?�0\9��)�L����a�[ɫj���H�`��>d�|,@�HU�KpB�O��1�(A���r	�e谖#���rt<Jv�$ؿP��d����u���n�B����L/�[����v�S
1t�;�����E�-	� ��6F6������B���A��!�}�huŜF��V��=���h�4�K���/�:��0��:r[< #�����s��a�'���X͕�X�)k7��ʘ�t�~�NRx��/��Z��d		�l�i[8�В�ZC���ښ0vυw���T��@��5}�֎v�@�3G7	��[��ũ5s:ሂ�=bf\dJ��:�4:e�ekL�z_����~1\5Ǫ>��N7�g(lا�v�&Ǖ��>,�d�۾T��1�l^�p�,�E�u�z�^�νՒl�J9�w��4hW`��$Fsx��	"o�\n�P��D�A1�B;1��������Y�kQ���,��/��u�[�ध�Ƕ�[�M�w*�]�E�-��"��X��:k%k1�/�sY��N��#n�1������7z��+���[j��h	lq�xvdO7jM���2����,�}��"F�و,U��ppo�]�G�[��h��tF/�"(B!� ���-�0m�� ;X�<o��5�Mf� *Q������i�`��"�\<�~B%1�g2lZ8{YJ�F�W�~�Q���$4�J��h1�#�����/�r�}�P�0R��OJH�� >���(������+��3u>j��8y}�oUH$��O��h'b������?��!���8b.;�̷�H';�9[��_�G��a�?�O!���+L�m�~b���n�)��ߵq��+��A)	7��ЗU���sn�5�f������lsIb���~�;0����)�z��jmU:t�}��ݷ�����:���Dt甴L)U�K����X�s��\����*9���u	0���Q�t$��j���"���n�a�'�μ����!=���Kr�.;� g�֟J��ٮ��T�-�b�$5��{g@rt�.v�^ہ������_SK!�3��-�Ƃ��%��Z���_�7��$� ��
���z��}r�&9~��q2��E��=<��JwT5�ۖ�K������zZA�p����9jP�NV]�c@�//ӮB���)]1�R�-M�֍Q3�<4�F~��:�|-`?�0���>1����p%T|��2ϕ>'#n���wqs�{���aZ�F�wt��� �����'�	��6��M��{�ZY���6	 ^�Xj���䖛z_�ٻ<!��eW������i�@�Q 3X�z�C�Om���OMƈ�"���4�I�.�����-|Qhnн<����h����v���S�xS-I��cf�]��(��̼�zW�L�ٓ�F ?���-�	⟒3E|jCb�~J-x�遦� ��ڰq?�e��5����z�[Z�Drkg���ԓ�}��	t#�hx7H���J���/��^��E ЩC�����F���7nTs�E9���X��a���� ��Z���I�!�y��bs�y.�����F�'��0����鸾����|�~�m#:�NstB�M�mu�]|����r@hO���$�%��m��>���=[<ǬPnsͯç��G��^�>�0��*���)t�eG��n�X ��xYĦD�P<�m��U�bBYݜ��/.t5���{=�)T[�[��-���+K�@z��� ���[��GR䢱��w�y��E�̗B����e8<<��-+#��3r%Ґd�c�����<h�������u���G@))+��GL��]ɹN�5!�4�tS��0އ��58T���<]��#��7����9n���7J0T��7�_�cL�P���Ђ)�WaZ���0�l��5�<B-6��!����F���.���Kr�w5>���o�Ph4�Xӧo�"[�Z�gg��F]i�R�	���a��8�?U��Sa��*�X�cx���Z���q"����wԁ���A��w#k�w��Z���H
�"f����$T{��$�%e� #Jމ>nX��x�(�����+��lؐC���ĥuݾW۫����,�cC��U��3pe_��δ��e�Ҫ��A�����s���?��bt�k�^X��V�������#�'�7�%���� e��ی�����[�.�����.�i�217�/�����$2<��΀���"�a��z�f�N��.���qvٹ�͋X�So�`_����K֩t9�F1#�ߛ���J\p��2��EjH�bc���_[f�Z-���;k�'6�Xr������C2`�0;N�eU�,waV#�����S�9����B:��vf��*1�4��܋��QNލ����V� ���LB;�#U���ۑ�3p(�{�ߏ]F��� �rlo	n��l�j���oSW�Y�ݓ�!�`��/d������4�u�=�@�9'�x��'��: ��A�O�Ҿ���l"��Oߞ�aX&�l���F!�H�~��r-L��s_#cZ�y!6�Jlq-�z����@H����/p��h6�Fe�"j��]�L�B���_��覼�!AQ�)�^"
A�Є@I�z�#�N�S���s5������A�V��Ú�#����B��+Ȣ��Q�T�Q�U���������_������m�iW�nYMv	<Ѕ�?��V�s^#!W��/cb���skggi(a���Pflg�F�?�t�B��!�:!��8����qʭ����\{ϵ�:�Ky��_C|�T%Ҙ�,i�^�����m:T��������b��L'	�J���Y��kŨ�[� ���	|B�yw����E�����P�޴=A5�BU�zH��m��t�E��fx�7t6SN�(�[���i>wY[�X# �s=M�����8�c3��_����i��rmbP|� v���7[��s)�cΎ:?�J���Ŗ�ғB�GU�I�?�9q��h%���3Zn�#��
�%��ʴ�>�-_ue%(긇J݀�,-�zӭ���4�n\��p����&�C�����̅�F����u�8�Ě$�7In�_�^#�����ب��l���˶�NR����`9�Qf�z�%��s�'ZQ����#]#�@,|�=�8F�lҍ�8�����A6�D������>�qY߮��+��;W2���6q�7�@)�,,6WdR5�Џ���k0��`5��3�^m)��#�����#�1�6�/�5J��˗�q�̡�'l�����抦�,�m����t��5~���)�(e�A���LE�R�����^����� �o<@y��iR���Z�a��X(�����(���̚�b
����X �OkO,�c�����GC��2�zr�>�GYA�,�(��Q*��f&u�)Hu˝{����a��ӷ�|�I�2E��y������YMV�"E���t�-:���-�� �#��lOOuq�N�Yĥ�6g.���[t�f�*-+��5>#��"��4�lNc�Q��X���]�V^K2�j�u�R�M��@�P���{���R��*m��{��	�ɫtC	Eϓ�������2��
JG3�p�����;�U��r�:8T��2$�]��������
	D�dS��K1>?3����+otG, H��Y=���i���`��?����D)F��E�y��4W�M��:��F>*�@���bʽ�b��)���[S���e�0@UŁ�u#�ʋD٥��"�d���~ˆ��BQ�K����} �xt(�ý7l�m�l�Z.�-��|�w&͏{�+�\#˯EfD�fJ�YC�?�0s[wT�?�Ix�E���?+x���X�}�.�S!K��5�֑�M�9��W�d��M�+Ih��h�H�9�4�[�k�0��٪�x�G�ȸٲ��m.�8%^�ѿ�R2~6H|��v�*'4d��~�i��Epv�'��ߗ"��f�?3�&Kx�a��D_�S<W�$��Z�`�l�lS�}�dae�QM��P�ۇ:ܣ���T�����]6z��<(q��"B�g|E��L��m���������ْe"??��F�k����W � &��k�H�ˢ�R���u-ȁlv��rO�J(J�Ɏs��jg�_�&f��IP����n�yf�=yMC��1¥��D��EP��νD�"2��Hj����5j���j Ʀ8�S/^�� �F�v����|+��#�?�~rc<�f.��67��A<Jg	����"x%���>�qG��+ֽ� ��&�)N�B�3m�Q@��'���rh�a���,f� k���Q0�A���5PC|����9��6�$��nѯ�0'd#�@a��ؿ�w�r��UZ�{T�!����YK�P,o�kԤf#:��W�㧢:�H�I�Ӫ�μ�?��CZ�F�r΄x;q+G�0fٞ0-zƷa�>@�P�J�Lդ��o<_��?_�-��c��r�����E�)����NF������!�%4���������8���8X��TKQ[���.<����G���Qv��~=�E����d�����S�����oEJj���<�)�"*T���_s��'���Je�&0��zt[�{�958������$T�8_-W�As-��ضY�Uu��_F��Z;��vi���r���������|W����k�w�O�%f������������&�����~�+��[(��d��n�rh^T������h�Wk�H
�ZK�*2y kZ�������A�6�͗�+{��+�7�<:RU�j�e��m���o���۩��+�}��`���%��:%�ߧ0`���{K,ʧS��Ϋ�S�~-5�]���A��Zp�	z~��f�|>ǽ�j�~.�=zk$���緄Qu�u�p�D�[nq����Y���"G��yI�@}Y�������9wS>H�=_3��f���>��]ȥ�йæ�R �}��8H��q;�B�d{c~��>v����㬚߶�[�D})!���0Ġ�dxM��]�E�鬫<�����`{H�?"n�P�,~��{�cٕ�N��q����Z\���E���V 8�C�V���C�[��{��^��8��Wňt� �2^�v`�0��
X���ÝT"�����C��;i�&G\��L:B�i���i� q�L,��A�8<�l��{!�Y��Y&�`Y�����ESn��Hx��)R[��w����>�y�����/6h��O���]�� �}�X��>���~p1E��#Փ�H�����
�5�q�"fM��,e�g���
�A>���Y���/��A�t�	{F��n'�U���?�,��{2J��.6{�Z~|�R����HOi�l=(:�^�O���k�K_����s��q�x��{��dEWC)�^]���^&Ђ��6BN���=P�I}��=�/w�N��O&T%�����XI�~nxm��l�ϭ�.-�a|�k� �5;��n%�̮e&'X�#^��X���D/s����(��G)/�I=�
E��U�ԙ�rNj��#9�G_�-Ra�g:0�pb�����
���*���9���1�z�����5�Z��+3zAA���'=3�lw#��Q��N����w<jV4^ll�o���J]ϓ�K�cI-a��J�0��+:]����,E3䢔��jq���� ��ɣ	h�������5�i�6z�	-	��Z��I�u^PYMҹ���k��"�R�Ys�Z{K<8{���;,�wL�߾)�B�e���ҥ����~��;lH���*����c��7����)��F�]�v��9�p�oC �[���7��^�g��Mg6�r¬$p�!:����gE�o�x��0�A3��!�m^���П#·%��R�^���%t��;��M}�N��X���� ~�S�J��� ʂ�,O�N�0j�T�Uh��2�)aRԵer��</%���#�d�J�}��r���Z���M�&�����v�J�������%	8�( �N�V؇a�xp����*[�r>=�og"[��&\\%����L��Vwi� �#@��>a��C��gBϫ��ЁJ7�xa7b:��*z��ܼ��L��C^�\��~�XWSK�Hcv�+���c��-���\m*x�q3�K�&1�Γ���^� �c�S���� GO-r��9���"*WN�7k��4��?�6� �!Vip|�/�DQٮ=tO5�nh0��eA��v�hg���کC%�[�T[\�������>�p��@��`a��oƄ���?V<CSA�lBQ���w��T�����<���\)�_�M�ïoW���LyG]b��_�J����b�RQ}�Ϧ<qĤ�rHR�v��%x�h���hj)�2�L�N�jΏ ]4�@�ז�*��~������z��!"�~_��>�?�K�In�G��j>��ttسk�;Y�U����o�3z�C�����+�^ԝ�SKl��"m,�W�]t	A>y�X�=AY�#JX��<~6�	������0���Ϸ��~��Ëפ��F��ꨓ�*�?s��YI���խ{��^�"��OSBs�PW#n�u0*��dQv�t��=gP�M��<Enx�5�����Ќ����yJ���m(Q�d+��G]��S�֙k�l*_��m�0�nbR�ܚ�M��ţ>��bV�63L�d�x��D|)�F��1gx^��m�mDri�n�a9��hG^b���fu�X�������kr�(Wa��Gx͢����M��|�5?��!�����E��s�y�a�ؚ�H����!��L�o�x���8�Y{ 4�}��G`������g\nLR{�7��g���:����/�����?q:�St�ү?M�`��w�^�F�ո�(P9A[�M\��#I��C`)�~+��(�ԝ�J�:Ȕ?������b����]�5#/\NZ\G��l�a5�ɽe�ʮz�iP8�U),Q�:p-�Z;����9��2�Ab��4}fP�
N��[GT�����]� �[Q�g��X�-��9
�%P-hi7ؗ�қ��1��ہ��vI;h��R%�G��ןΫA�Ƨ��X�c#���+��N?��;כ�Y�� 9ɪ�.�
�"ӫsk��N��L@��\
��N�z �xݷ̭3����"�̆�������y�0����5d�UA���]I��8�$�R��P%���%�*�`�#��yz���w�u��� h=��0�W����,�,��m���v�VX/$���7��e�J9L2��`a���á�>��Nh�����o�1Đd��pB�o�KgkM���ㆱ�8^�[��l��Z�T[j��[?��<��([���iQ�W ���Q5�K����e1��ɋ�k�0�lL���6׎�Ю4�P��)[-<�K������=82�� �o%F^5N�"��Τ�|DO8���17���xgs^��	���w	"�\I�`����'`�w�W�Jj�v ��颤 �|�]�¦M�٭�R\+TD)?͎q]�T*'�Z��ڥ_D)�BjO~n$����gf��3�C�ۏ�w���H|�Z�z���&ꩻ̄LFc�1b��8����A��J����/A��Phe���,'jA��?��"x��+E4Fq��j㵑����(�j��^�Щ�gX{J��e78w�fu�7�����{w�%r�;��닻">S�n�\�cel�"�8F�_�#�L<C>��w3.��g`(���fjmC��W��������خ[��h�H]�.>hɁ�ȧ�&L)�� )���ڽXG��Ϲ�	(��;��%��E��;&�*�fYv]Y\*&M��\%{�~�Uz/�͙�!)���B�8!�x:p�'��sD�!�o���Bn4R������.�cC?@E�
"P.�ul��_��^
أU�Z�7���3P���]�����D�4FbaV;��V�7D��دC�8��S�V#��@U>�i�m���6Z(X��h��I=m^�~u,���S�U�s:r`�`����p�⾩�̗O����܆C�Cl��n��Ht٥�S���o�ā�f
-�}y�������5 Qyw+��[�@�ik<p�=��Ku��M��=(��ǻ"[��!��*���a�C�d�,� ���wc����������1��"8�/C`�[������ƋW�>4 ���Wk�fK��֯,xcA6����e
̯��A�D�ҶU/�ra|"s_V�[�|tտ�X^��e�sV�ٌ�^�:S{��%����+NB������R�S�.�bL�E�q%u:ٌwG2�G+j~Ŵ�r��4e�E,;S`إT[�d�_�Y*!���k�P�� �W#��w��e8M������y��'�UgW�^J�8�˴.Xў�Y�>t8��5�K���u����U�P���ss~ʍ�T5IyP�x[����4�'8?�R �
���7�i"EM�݆��]�<�����%�B���S� [�Mcx�� 𰷰�ڜ��e��ߛok�ơh0��c20��(���qQ�,��n�����vxP��%��<�Qoғ������9��r�%I��Z>J���<\�	��J��<�	�̂Ee���{����ˊd~����LlZ�jpaq�z�W(�����x�;d��j���I�V��x����o��S������Nl��G7�^���n�I-&y�Qf
�Y�g�p 6�E�f��˄���+�P��L�8h��`�5�	�$wy�7��%����=E��K,���XPyb�Ţt�x�t�F�l�i��m��C��;�����F�)����C�_�ƩާW����bc�D�\߅��v46����˛��y�N�L��b��gןP/1r�3�3N�������g�7�Q���t���w����:K�EbL>@�`���]T{@}!�-�q�Pz]?B�{��b��������C�88X���eE�Öܱ{k��W�z�fc������2�.l�8���yB"?�����ai� �hy�����hb�ԗ�����z���k���ؙR�X�����3�%�x��m΅4�����`����ì5����V�?���I������P���D@Eq�U�D�~�?���͏1��y�<,���0ܱ>���x��oL��ii��Y��$F��*1.z���I,��ĝ>4* ze�1��Q���[������VBK0�7?�m��![��-U��X�#V��5Ļ �Ϙ[ݩ`O����Ù8�T\J���a'�1�S������|�JS���i��D�D(�]ԉ���1idf��m�U���f�}K��ι�/i_�KV�~�1��D�{�3�Tdr������}��늹�3�e���9.a�'b���#,��A�q��w�	�A���z�0oVX�z7���A(��/�c�4�ْ����;�dz�J��G�k`k��@*$����۝�Do\�ř�)����c�S��R*��}�Q�,�;��5����B��X6:$���D�ǈ^K\D�jI�G3���5"L��l�U_��͟�g<�xt2F5�o��m�zF��X�p��j2�'�l�K���,������[��� ��ռ�!;����1�����UF�I��"}/���s��V ]��Î����>{5%I*RI�{�7�1Z�̠��&�~�{0�)��/Mz�G��<62��Q�%�g
ٗ@�]j��:/��e�����q[����
�N[Pŉ̴�E������/��-���ٿ(���k�u� �\\�u��zK���|�Q��	�<���<u�?4s3C�;e1�0ԟ���T`��Pߧw@�cqp����cˏ��_�m�Q;�g0�%���U��%�pva��1��p���}}���7��5�r���M���X�7�O�!��%w&����P+��M�a�R"��{�T��[3�Fm�[%�H��ߴ�s���<��ݷ��ξm����#���P.�f�!xM�!����9�b���)�èM�;���z��ra�<��
��m�+=�@�͞��Tw��3�9�'��ft�j����R[o̽�VH@~/@��њ����{FW[S(�s7��%��ϓ#9�'�ע���h��"���vOBA��*���h���/�ct,�H>����0�B�=!��9Y
_�5 ������O�"$��gb[��m��} 7���<&�uxV(JO��/ɫsj�	�2�����ދ����p-�>���P��|�vk�(��V��T�lB��
�;C��fC�ʛƼ�x��c�Ùlh��,��6W��9T3�ʏw�Ikl��{S�P�𜂓��/�q�O�؊��	jҷ�y^�	e��*ǒr���'?�b,��@��a}�z�}�D�v�*s��r	d!7Y)��MK@9���h�I{�����W?�dLd.]	jj��kz�ьw�9�5{����U��p��Ϸ�=�HP�mh��Rs|��s{�O���ݫ
$����-%����"�i@�H���[3�RV����A��S�J�)���k��ʮ��z&�G*�SƂjTJ>�T�'����Ҡ �����B��D�/��dCF�����=>��Oa򂏥��Z��n�J�R.j9��Lv�Y�}&�`N�7��j?#,)��OQ�gda��6* � n�IфF0Χa>���%��D��ȶ��afj�D�(���A���hq�͉S�Z��zwKe$y����$�37�Q��X�1�Q๢1��nq�B gݬE=���Vn����%"r~�T߃ۭv&�f�����^[�4ZZ"���Eİ�s8�|�|~���1]��\��rhP�n$t�Ы����LR��mS	�Z���QmwhK���{�ܥf,��kp0U"�Y��\设�o�kW��0�W����bu'�� P#���a�so���C�Q
�h��Z��/�TC�>��>A}���a۫�(�.;��	�x���K�;���?�^^7��3��7�ҧjKN�}[�}>��@�J°<m)sC�⏘S��c����G3臰eͻ���D���TA�a1����!:����������W]@|��ǥ�Z����~uR9�}���B��UFvkU�$��[��Q	����I���{��?mM,����8����ɮ��Q��_�e�n!1���ԇ7yz�&Ю��/�*��dǅ�M�A�Ɋ-�>�J����b��y�[�ͷS ��k��q����T<�}vѸj�Mhvٹ/y��&��RN�jؗ��>��ep�跞��t��'<ҟ�"��滂1�
�uA�=�M�'�@kn����w�3ȉ#<BV��?_�p=J(���MIQ�c��C�slX���8H���p�Έ�L�#�N�%���9	�:mR�Fh�o�`Ӂl ��<i7�X�U>���Q���p+P#"�@��93*��U3�X��� a��'?V����3�	��"]y��g�QT�;��ө-�� Z�q�k���d�@0ݸ���.sJ~��v��.�ᝫ/���F"�eš��Z<&Ħ�������;A-XYF�Q�V_uS���A��ɟ�/���?j(�K�('f��vA��t���:M����s-�{�)�ّ�a��;��y�<ץ�D	3��a��u���{j%(ޡ)����Q��L��(���k�jS�ʖŁ�d>�T���vH2h=���,��Þ����uD�!2�[�7Qc��?�ՑrCLMn'X8T�ߝ�e�,r���6��^] M�j(�m�m./�|D��)�f!}e��Xl:F}�i�k�$��˧IH������s�EA.�D4�D��i�(�x_�E�,_�4�x�r�F�xL���g�q����L�Rp�p�|��;�A��	��5n��	��jğ�c4&���t�����@&m�v��O(A�u=(�ou�����wZ�=�	Ef�W�i{gA<�ۧ���)9�����d�k+Tːj���}=���~��@.�	�L�nsE(�ڝ�f{������ ��W��Ku�s�}�;$������K�wsդ��7T�W�����$e&�Rv�J��J��'��G�w箦H��Dk�0M�- �����\�I�$ ���i��膜��r��h���C!�����6O.n��`��$M�ܱ&��9��#�C���>����C�d`>ZCpd>��Z���1���޾����c����oٔ1␄E� �ұ+�+	1�M�my0+YhT���Ev��P�࠱��<�'3,9�h�/��~���p0ː�]W_$�*�U�m��F}�A0 ���th��@	�������ͦ��rQ4}�v}���w�Ĕ�"�X��#�@��FS�|����� ^t�Y���Y>Ψ\�7���R{�8L%����̺Qv����L$�aT��*��h(�)2�r����ʲI��oX%������Gd95ߤ�Y�Ӓ�(��06������Y���;���Bk��Q�pv�}��ri�6��f[�ZS�f�L GHm�?���� �����nt���W���"�Z<���/]�CF�0��V�o���DҠ���I0�X�����f-�%l���'����e�T6ф��#v[h���;?��ABk�av��	ߡ����)�]�ᆡ-$��u�gb����=Lp�x���h����HB��Ig�ڗQ���������G��F��4���y��%�6�ѫSm��DO�����>LH/�<k��^|1tV2�7	����&�;�c��D >��Js�¸d����;|_���u�Rԏ"O9/�����և_�x?��R��|	�A�@�g�Ed���2VBHۇ��2߬��1kQ�\�7�8C�ϨR�?/��)��o�ž�O��f-z��AO�R���F�e<�Q<�u���zn��I��ѵ$)]�<�/�'��Q�\U�5C�<y;!�Ko�L�yR�O�,���
�|ZK3]��J�l!-Y��)?�����x�~�MrxRX�=�d��r��pU�d+���[:��R�1�bf�$yT�d¯��0-�zgZ�]`f��,Iҽۀ���g����1�E��֜)�8��R�e��殛'�ZQN��'��{h*��0�����[��uam�	i��(�Y�M�o�5վF��h�8n�K׿�}v�#��+�S�p����!R.�����CM�z�l�æ���v���~��S<Qu���$�$���GT�q�r�͐��~Y�9�9��Y@�8v�V�N��R3PU��æc����X�H��@w3=e�&,�7��+� {0Q4��e�J'
JT_�$1�}�=S{[㮵�P���ɸT5(;���?��×�(t�h�@����U��^լ|���\v.Gj~
�`�����=�Ii�͝+�e���tP�1 Ph��m��ji_HZURz+-��z�Ƶ�|����.G0{,Rt���:l
Ù���+�k˻��~B��ј��	M1��x=*� 0���U<���������Ӏ�l�;���5�����L۱X$�!������޽-ˁ�PU�ncx^�-���@ 8��e�4`� ���~4��A���9/v9���y'.�zw����s�FE�>8���g�t���P�+�#q�K~NM�<�����*l��P*V�ZL��"i�͇BI���c�j���by�m�(P��z6�&�a1��z��X�m����e��=;uh&~x[�%�殯�����K�ډa_Ru�#_k/u���G�>]g�` D��Y�>-gaƙL�-X}��I,��q4O5R�]^dkE��u@ ��o(��s��+#�m�PCK�@9i�N.R��!wH��ӢΝ�"}��N�~�l�Ȁ��e"�S 1͗Փ�m�Y�q^g]���
��B���r�����<D=&I��\��t'����$�Qɭr�]1�殣m�IN/��Y���{x��o��v<O�0Mr�'o�9��OH�Y&����{_��VT�cz���t��	�3P��%�_��eLj�]׻]�Y.<̤�����KqZ
�a�e�"'�����Վ�5E�.3| �Xz��:{�8Xbq"�Ό8�8_��Ll����b��J�����L¨�qLk,A}�G6�؀ժI��{*owR��A�A&T���3�Ԫm�j\mof��J����I����ŧ_;F�2�
�����]��'�Ck�u�:�-}�~c�-[�x��1ٓ~���7�3�(��c�߼�Pj��ݐ��1)�Gٚ?��R��ؗ���'h��Q|0Ϥ>Ϋ���sS���/Om��[m����q�?d�JK4��m��g;>K���"���a�(�.F�B��ߊ�)
Q�'�o��߹�q�_��+�NN�w7�x� h�g�G~��!�].�0�%eKt~Ğ��Y��*��7�?�`VZ�*��L��� �����
�ɬ�W� Β(u��6-8^A_�IoY�8�ݾIoށ$�`��?f:��1��9�t��k@u��]f�JT+�p!��O���L6��'D�Wt^-�jD5��Ltu�I� ��VrJD�F�>��f[�������4B�~ˑ���c%��,�%9��p�G$3w�R��T �$%�!ce`mKz�W�n���5�'�
	�SV��g5��y9�5?PTz�؟�~1	聾��uh����W�����H�u�����Q��T_n�(��%P$�U��k���?�p�'�/TpX��ĸ�N�<�%���Q�� ���A��t�rQ\�5U#�-x�� ������Uޱ�s�i�������s�/{N.�$�{)*��6�Ūl�14_7T�U�	��D��D��R�;o�d&i��(?^�����@*�����C"��P�t�@��Xl|��
s���|x�s���&\H%Ԯ���&�nVw ��5��H�伿I1�d�l���q��۰JqZ���'��gZ�هc�'2lZ�$s���_pG����0�X����:���G��8�����t�s���2{v�:��Q�q���y	��c��D���g��kR)-��dV�����i�/I��/�e�b�4:����'���Φ�EG}���;˘�3���v* t��(��GJ,6EP�0H�_�x��iQK���������ġ�e�C'c���F�50���pB�YY4�1��bU�zMz�g})�(, ��D-��q��H�7��41�q#`��'(V�]�S����q*5�y�"5uG�o�}(����Rs����[����^~�:K�V�y��ɓbG��6qԛ�g ��_����yx�6��G«���0��=Ѧ�&y֐���uEm�7���*k(
�����B�6�]�6�������y4Y]�j��z",Ú�3[Or$N���hMJ�ɮ5���sB
Z�#���:sx���xV0�+Jq�{c�xl�^$/����^qMf����\P���r�z�,�w�$ƅ�{DP���1%���1�����W�� ̅e��SX>���ӿD�؇|,J�ڋf�yO�a��e���-~��`v���de�[E�t"1[�B�)]࣐�Ѻ3lJ���T�!P:�5Q4O���R>5yGڙ�O9�Z�75��T�����"�<���:i�yo�W�Ϸ�
m�ʡ��S�5�X"B	�V/1E��㫬:��e,����{#�~t[������"�P���P{������V=CU��W��� ~їVO�ɤO2;}V/2!�ݓ���RC����I��s�7D��������O�D����j��r[qM\���u)�R���N�J��Q�IE��m�1C>�m�6�Y3�/ηT�2�5���T"�r�2�}����4�;bqH:�XıX�.L�.��������)�����71?ȓJ������pz�w�L�ڎc������vw��kn���(ٕks�
Ƨ0t�O��\���i�H��Ŗ��Ѕ�_#Z�b�dX 1�}�k��`��l.U��Ap2s�0����~��<p>Ƨ{X�K�Os����/3'AW~�3��!�u1��%.XL)�ݗ^a��Q *L>[����n�i>��ǫ7�I���G��Lf@�O{v�Ծaȭt~�	i�i�TӘFeZe��9`��$��Y�������:O�-m;8�x�ca��.��d�GC���/���@��&@��i�w7�7��k�Te0>�Т��p���$� �3;�i�Y��
a�_`|���WkuK	 �k�����;������Z����v&�؟��ܠD��޸�5B��Nx�T�lb�9*[�(���+j�]��9���ZV�-S{��-��
�<��P{��wꑊOfasq+�*�c��l?��0�Z!���^�zXh�z��z�v咊ٳAp^�x��5��ll:�L3���.ƾB�ז�2����`�g�6��V�D��s���\�d�r���_��=��96����W�:s����9�p�R�G�O��j�X!'�_Z�=]C��1�"�t�*U0���'�!��s���$�h�RL�M	��Hh��h����<��~i Z��B��B�X���t������/����u�yn�i�28 ��.��S`0%ɮ���]�����#����^����/x#�=:��$�����w�/�����v�ΐ<��qE�
8������̅_Zp��݌�
eG}E���������*�%�&ur�m�k�Ci���q��
8c�c>|��1�S#j*@�%';�dA��+E:H	�iN����`��q��m���|���h�Nn=A���R�9�$r�(��2��~OXy%<+hz�����`t�ή_3�R�^ sCI����TX0��&��]$������<eY_[� ̩Χ��%Y�2W��D+�VBM�1��8�y�b�Ҁ��^�NhV�]��A0�kW��
_���W�����$z6?5Zc�U~�|E���Y�Igǅ��.<p
�9�殢}#n����Q$b՘�E��r��K+�]���!��ꮞō��ԡ���	�#���I� ���ʘkMH�s	�ۙ�T�&$���L�3'�+���أ�>.фS���e���R�Me&@7Β=��T�Oa�����CĜ���2���J����^�7��kP���#���8���a/r9�"rup�)�Z{&��m��ċ,�� ��<�s������ɯa�����z!�G���ˌ5�z(�58��U�����%�z����p��岔	@axp�z�b!pzb�:.���x���6�������aG����,Й��n?9U��rLR	cq�Y֕|f��3&�Ɣt�<a黐,���4�+3O�<��۞v�p����|�
bg�W��yN-UN��N��l�b7!&�*ڬ�ؔ��c�e[c�7$�OP@ۃ��@���#�,i��G�G{�u`W(��5(L�6���?��y��hq�06w.ԶŲg����x��ܠU5�?.J*��j,�2Sg�*�t�~�J��Y��tE��af� 3���9�a���nJ#3)�8R�T�Ș�
tM�G��	��~��uI�,�xh���Pr���U�a�^�af����[���o�ٺ�|R�E!yI��P�
>� ����Ƹ$�|�o��)0�󖏄ëC�A�r���<��@��cǣ2*k�u	]�i�
O@\ۉJ���	�����!�6�i�H���oC	��v����so-�o�E��`jc)�hF�Ϋl�� .�eܞ8�����q�m6>c��ON�"�!v�3�[l����S#%Bt��v�atn�xt�<�C��Y��l�dL�A��(�x�&��4�����G	�i ��M������_��]��ˠ���)Y�~���k&HElsGĝq�Tх����4m���W�d� $7ëWG�jǺ����I*�o��7�����`Ze�!��&$���������9G�]`�\a{�� 
qjԪ�J��>\�u��hё1W�?
������������=�3�W���~���z��u��#kF�pw�U���$-e"/V��"���]��U�����H�n�V�W{^*�_�W+,���u�`7[�����%���!�Ռǎ���hzH�@ؿ�E��(fp(8�|zi��waΣ���b�&܊�'�X��FK�����Q+b^8���HG�R�g�f�*b�@_�o�+�֜��k)X��sC$��vC٦���L|�5����i��l�(Ȳ�w�E����/�w'�Ӽ-�%�E���PDs�9=!ܥ������c���%�-G��.��q��R�ԛp��P��Bo��'�^���M��T�տ��֠o�3]�	����w�Q�ƒ�ȷ�|�P?<���_�Ҝ��$�y\{��.�V��̈�f}>maO/�#��j]C�8���sqE*��mb�n�y�ŗ�\��ܷ���W���-�'{`�����4ΰb����ŝ�G�aC���ک�ӯFR�	��8�U�>�`?�K^��|I�D� ��ʇ��K(��[eOA��n=�mJ�PLu%�ӎ�R�#��Q���a�M�4����U""G���u��ς�<�lh^�^bf��4lg��M�~�4�\��ҧ�B�1)1R�XoD�g��>Z던H�V ��pA��hTA�ܒ`y�JOJME��������Wk�@<!��r���.�0���xl���%0��Ȋ�Eu����eD����l^I����I�3��:���&f�~�<���YZA��b��ٶ�!�%�OD$�3+r����joj�v�6��@U �V,���� �Ȯ��K"�1����AB}BNaJ���In�
�[��G�1�q?�?�;6�E����\YB���j�|��=k�E!Yb"2)���F�*k�{@ �[%Ӝ�Ea�~�f�2[B��v��Ԗaڅ"A!+���W�Ҥ����,p�l��v�x!
x��и�����7f�a���C<<���+�=S��#&t�� �s��^լ�����F{yx Q��ݔ�5!�?��6fKA�.E����|/��
�ֱ�1<Z2	js_��<����^��	oiȈ#~�ȃ�eUP��Q،1F��G]45��GI��ׇ2���y��n�d�!,���S��̤�q[�U����ۭ$��+���[��]�:a\��z<<R<Oh�m>�}n*ƾ-'zv\F��I�n��/�T²�f�V��m���,�K���@�=8��X�Ef��e�b���_���)�,�C-n�X���5��>��#���|�����l:VK�N�����E�=	,�=%���#U��J�_uY2]>�P!<b���3"����Ƴ �:�Xͱ���\�!1l��a����������#3u��$m�q�J���{Z��� ޝ��{�H�r6t
r�MW=@<�5��1�y�C�8���D�V�c�e��C�����B��+	���q���'V�L��"���:fA�yF�{��Er\o 0ɒ���&Z9mj�^F���{���T<�|-����|@;��s
��u����ߨ<�Ry�6�N����9Tw^��R @�2&0��Y�鸯O��#0i�.�$��P�te����7�q�o�X���B�jis#Y��^��ə=	J�vM�Xor:���z"�8v��B�9mi�K��E/f���'��R� |;䒏��4��Y����!�F��q�����$?!5�S�ے����H��YC�Z=��o3҉�]�Qe���-�E�a��y��n�p�C�}Ȋ�5<4��;B�'�\��˔![�l�����g,m����)D�d{���^�i+�h���E�[j��g	�lR=����4���7P*n�m�,0;��#x�i�=)	�-��>(�Se� ��ݪ״U��A��]�ov�����a�q�i��D�wF���vR��kU
��͹q���E,���[7���3ʔ�䑊��e&bSw��d��#����xE>�t����
���t0UT�h�?�#z��}k3G?���Z��Yrhf[ZѬ��N�*'j#�0��ž:4�~��3���~1�#��D�i���-HP�1�]���m|
tG<#��\~2Ӿ
J�ܙ�B�()�j����HP$zkq���4�Z"�74�Q7��Z����$N\bԺ���R,���&����Q�2�o��^�y��1̰����'2�T9�����po�����ii������Q]��Tp"�cZ�.J�c[[�#��;׊�J��-7B����d¸LfHy�Y���.�1��ii�-8�m~Q�DQpq�P�88<a�d����>�EA�b�тR��c\<�:���JQ!�>G\�y6J���L�����4\��$�	��S���7u����l��(b�_~ë�'
W[n6p�"�ˑ���mԻ�ԟ�P���g���17��1���(I�m�l���6�]v҂	`<t�8���v0$�Q���ض����Q1�BR �\U|,4�C�˦�(�>O8���V�5�3��%�����r� r��ϻ%5��9����*���3���IXfF�Q.Iq[�h��4�?�x��83��5$���i�jհ�7��KA7��!�^O��b������ܣ�%Ĝ�3�O���T0NoĺGت�$������xC�hi>w�8����č����+d}sJϚt�A�7��_w�..�xAu�*(F�v�����D��nb��g�i���w7�����V�-�ur0�Fd�����5Po&(���G��ʷ�=�L(љzM?�X7��<ٹ��sLj'ّ߬[�j�k=9�A��z��e��?�!�<u��Դy�7���4��u1��X�>�3&�1�z����D�ǎ�jlB�6{�؜oj����։�W��Gd\?1�lӸ�,3��÷�P�˱�8ҡ#d��)8�8�[ˈ�;yRꤐ���w�T)��M��CmnfɈh�cJq����|�I��ǤzʉǂC;W\(��7��p�������UT��ed#+���q��F���Pft���ᕽ��I.������s??�v{���V3���g-�N:\O�vx�[V�vP��%��p�y�1#d�pa� ���d$���s�����!<��v<�V4^��&E����/Z(�WD�/���o  o��;)�qc��9���k�ϥ%��w#U*�p8{�7�{�B��
�ĩ3VO�1�3`�p�����5a���_�o��T�� �l�������[~D\q �����%������94��G���֝�͡5�Qr�͇�؄:>/M@w� k��M�*��M�� �(L�0�:D��l�F���������	����J�&�cMC��e��#��p���ix�v6wW�ʿ��ݛA�E�KT��ȅ�	�F���G�_t��c�YWI�l{5�J_S`YC��.?�2�y�s�]�Pn{B�4��D,k ����Q���Y�cFv�����(���h8%�]M�R龧��ٸ�wF���Z5R�`�{�1F^@myp󝔑>py'_���"j��n�
^5\͢��-\s12�ښK�E_ˊ*��3�I��	��8Aq�9\�I/Z5�KS	h�{3��x{�=��4Uq���/����Eđ5�Ek8.[}�+- �!�F:�E�`D�;� ���)�Y<+h���l�3!���dO�`*�T������2&Y��y=D�4A��:l� Z?�7���F2�S�������5�gy��_�x}Qԓ�s��`E��X�/��V���Ө!9�tU+�'��({����B`
��hUc�2��A"���V�CR������ƉL+�
�s$�cY����tA�zWc�ҺJ�A
��SM��p���g	�ͺ�x��t3#-�c�B$�K��#l���4�)�A��7�]N��׹�C/B��~��C@��v�0+د�H��V�%Q�t1��&<�I�0�-m���$0��XL��s���g!�~я(9���_���,Fׂc�bDV8�j3:�rZ��*%Esi3mS�#��)�e��It��<�=�P	��P�'�[�)	�\}R����(���&�]8�\
p���8{���uC�EUW��P�-��%�Ž�-<�6��-�W�L��zV�!����c&L]�%wn���,�3��j�>1��Uu���^��1�Vk�6��>�!�^Ծ4w,JF19�!x�%.&\����I�.��G)TmC>&^�K
x����UΫ9𿽟R����[`���8���@B��%.��~�MRO�%	���t	>W�I�#<��]/�u?�*�V}5���"��.��tb�S�>Y�x�״TK�s�;��V%jq`T�W��d��b�v6��(glt0KL�����������B��*����k�.�&O�zo^�!�%��&(R��_���y~ ��
5���|��p���y��x��.��Zc7�t���tfL��-�c�ZH���
��j���:Sh���P]�υ�v��w��>F�`�%��M=�t���8�ѷM�P�$U��.o�f�:�h]��P���d&C�|v``�0?�p �`��m��2������FǬ84�l�)�:�+��,S�H�O+Q6,�jv�Rh�1��ұ�"~����&F@�(��K7�<����~�66�-nH�A��������Hh���p��L`3�}Xn�ߟ/��|� Ó��!����Ņ�`]�>�G�0;k�M>�������:�� ���1+.G*�^T�JeH�>!gJ�1J[�|S�^�Cx9�a��xe��|� ��NR��ї��Hr��������	�)�����}�`G �<��]�2h�Sd�1�d�)B0�8�&�6;Ģ�񇯌�%7zP�����u�4��:���|P�{B��h��*�7?�mR�QdCTߕbn���nX#���O���U��({��t&^*��H@딾����NMV��t�,���C@7n�}eNy�����+��ka�91����4��?�E�%��F2&	z�h�>}��-z�p˷�d�q�ąڞR�B�gm��r<��=����W	��T�|���H5��jQ�,���G�)��d wИQn�M�e���^�M�s������vSBwĢ1Ƚ�A��I����w|���������IPE\�:d��6��,�U�$t>g�\g�q��$LM�-|������-L@U��JE�]Z���w��8>i�P��hHI��4yV��V���؝d6u�WX��RGfUH$�\�v�N�JA
�7����vD����M�qz��)�d澋�e^N@@�
	�?.?�b�!�H?��gN.�l�

痛��:����礿�4��B��j����}3�4�P;(�9�:Y��,���$-&n�O�S�m�4?��U�?�h��v��'�!*Vz�u�H�<���y}��e@���|�A�_4.;�տ9aI;O[9C�"����$�♐��}dx��nsx�HV���}��O{+Z�t6'H�`g�Vh6�R����xyDh��3��(�]��y��rP����J�j��ϭ�EԖM�:q�.D�"�?������7��w�������ո�Q���qrLS��c}����������^�^=k��|�c������1��ɗ�s4*��l$Q���$I� �@�R�2�c(�Kl�RCb�%�FÈ��ֆ����q��T�v�����w!�k~�`�W��T؏�x�z�Q=�L�?zo�_[�Y�O��*@��ҏ�J����I.<�k!a�ہ�'�NUW���P�k�IyΖ�k���Ŗ����;�~�`�}�O���܆�Ɉu3vJ?�!����%kDN��L7Ԧ�	O�ܙ�?l������B���zʀ�k�N�yҨ����wc"^�@^�M��\̠)�|F|�<�0&o���Xת30�5����wl�ƹ^"�8�/*8��R�D�k*���g���.��wU>�=�Mgz�G���B��$Y��@j6��o&"5����"倗�/z� um�
��n���+9��]��g�~qس���R�x$e����
qF\]86��%s+/��M��+]�]�J���!��xi�-���[ ��h�;��'���NOa��C�����:�$S��#M�m]\�̃i�����H*iN�i��B0C�G-��Q��G�����K$�|tg򬩀�/SK^�5��42ٱ�3��dMAIq�J�!��->�jۣl0�!��@�?6�YZ4�<�RWp[���î}1Q�\  �>3���L�d��X�܄-,TלN����p�iO[ğ�Ʋ/z�܃�NbV�d�� �1�ܕ>��<�!�nr
_i���/���r�m�c��t�ιz���1��hQ�P�+�z�"[|��عf=���AF,w�PG��;%�X����Ko=^m��g\#|��.^l�3y�*:Wqc/�R9G�ͮ\���K�e����f���r�r��&���h2��9#I�m^q^����̛�޼�}gx+�n#"���I��X���p��O{׌��ڃ���C��ɯ�Y�e�\T�������gye#�1ɉ�W� �-�l�0�#Y��3/#�>�R3��Ũ�w�u�XX�;k��{���(�G<��g��UX/��?���T`���[`G�J(�Vx���/W�v�N*�� dx�����������^t�Ym�mQ5���-�oU"r�u����u��"���V[��m�<�E�- @���&����~���,<�8V����T��~-�G8�E@3Jڡ�~����W0��*�
�,G��{�"��-ȹ�$��{�?;Pv��*a�XѮ>d�>�z͌���M_v>���F�ʂ�Ӥ:zY��m���'��Q-Q�^c�W����]��5Zmbî�W����t$$ǆ����gPx�~B�$��I��ЍX��[���L�o�d�P1|3 I�Lx�����Ԛ����TH:8�S�A�fz�-7��[LK�B�k�����z:�*�i�N�E_E�s�4��=?�#�oAr�?#���̼��<N�^���s�f+���-X{:b�E���C���鞐"lk99�{3�M��ZRm]]�Gs�|�b`��sl������i��d]��E��'n��g�d��3��?�ɫ��� ����q���mB��&�J��4E������'��%���~���������B�
�M�sG�j��끿Y#K���@/~��)Cn�w{8�(�T�S@�k{{Ր(����Z94y�W���<�#��r@	��e��ظ��Ǜ���zY����z�׫.!�d	lsu���(�JP��0�{����&6�'��u����_�7xa����,@u���Mw��׌cz��w��Ed�\��Z��R����E��4��ԉE���d�v��Fs�"���֠$G�}�o��i�`9CZ����2�!��'�J��ia1%�����4J���n�+m�dG9�c���a$e��;��jf�%=t�@4?��=�V��J��{N<���t,�E�E^�q�q�yDD�ќ���?�n�$��Y�'��.|�L�	��Wq0����5�t�T�mmJOѕ���>�T�:�A�Z���z�4u�M�i�m?��':�1K]�d�����/���s��2�?��πKu�;d����m޿4�A��U��J/M���˭�%{�N�z}�qߪ������[�j�=�K0Qk<0����g�K��<�Af(��\�c�Û0��m��ڤt����Ǭ�phbn�u�6�c���A�q��-�����KK�<��:}D$2	��d*�.��w�zz(����+�u�*��H`|�O��F*C:S!���V7�/v��`��WnHO�;&�j�n�o�x(s�J���r��/2��v�Tj�,q���l��ŵ_!���+�(k�#*�2�_���<0H�:F��ƞ��CL�^�Qsr����#?�,?+x1_�y|LCL�L5q�����X�5p�.�d�V�p��f�p����Ƽ@�X&Y�����Ìʭ%��=&��U�MKD���+38P�ﹲ�H"���<��?g��p��(�>�1�	P昙��b����@+������V��t�nA��!"����(��n�;o���ER'M�`�]V��,K� D]>:�{c�I��Ry��"S�0S���i����vZ膷�\�17��If���qe���-t���Uq^4��"�<�/�tB{|V��#�\a4�VI���,���R�r��>B��5Mm�OGX�����:4Eb�"�l�!�ň��b��|�[2Yg%�wX.��7���yb��T��tB1�;Ӕy�j���	B�ឈh�Qx���'�Ԅ6�v��	��f�࢙@r�����D���*$S�m:�ٮЭޟ!�\C:@y;��lOnG:#Y�{jI��Mh;`Z�<�Ǯ�]�mM��}�k�"�����_>��bb������e�܊�в��	���b
��8�r�Lfv���	�O\)�$��Y�!�#5��=ա��D��x0+B�N'���_���P�3�HW\�7�U��6�ԎF�0�q������E��;³�J� U�h�c�vA�+Bt�;e�x��z���"Z젰�9ޗ�%.�qW|;��M�89?or��V�1;%[�T^�a�|��OY{���=ςX����\�P��5Uh��uvG�_�.1x�㊆�B}��.]��v�Ϊh�څx�QE�kпH����.gm�Oq���������5r\ ۋZf�T����n�T�uEo�u��&�lq;�r�]���J�
�+�M�6��̶i��`����s�N5��T�1��"�Q��!f>�]봰�s~�����Z��΄���i/�����1���{C�4er�1[����\mlE�I���P���zc��"��%��3�ܓN,2��������:L�� �B��-zJ�W"�;:V҇���y}�Q��_���UB�ynYn���B����_�q�4����SO�,�yX��9�����Ǩ悲2��������	SVo"�|�},�y��Ԃ���VJk���r�V�31�#]�&1u�X`����E.�n���w2?G�c�JZ��2�
7wl~�?�p]|,�&�m�)%O�S��=x����V�>� ԥ��;�W�t�$i4|�� [|TF�ۢ/R���Y0W��O\l�-��.p��x^��	GҡҷM�j���gE?O���s"��N:PO�(�=׾���ꪤ����P������5J�ߣV�A�(�؍M�z�}�<���M0' ��)6W5S��@���#{�2�q)�Ș(��gg�d��2�+�.e_)�YJ��ql_�T�_cÞ\f:��\qav�/i�j?��X����N�ԃ��`��)h����x$�³���Q��q����<��O�wP%Pe<Ỽ�1�}�j�9�D,���#���`6C�gZ���b�G3Ь!F�WT6ӌP��-2�hrI��ejcnm����^�5Q�rq���sHh�^�O�%��ϻ��{�Ts��,q��k���"_,H&7�:������0���^<}q�M�M� =9�E|Qc�R��(�w>�xؔc��l��b ζ-0iG��N�ep}�߾��.�J�gܫBxvܫ�&�`:���� ��4�Ve���v�T]��J\��O����r��Gd����u�n����-��l��l�j�D"����>D��|�!S���gH�/~�W� u�}B8K�ęd2���Z{�5	*��sO+�F E�W�E&�t/9�G떌�=J�ܱ�^lD��){�m4�1��';���VɃc�Eɲ��x#
���(��C�� y�J����C�;�G�6� �KC;��H7�A�J�+L���$�0���/�b��e���=�t�|~E��K2)nc���*�=Kß���훊M�8��uV�ˁlsPo��u Ў���ξ���;������'X D����3�ݪ��=ܾ0nH�j)r�ִ��iSͰ0�!��5�3g9��VH��*RN��%QD~3��=�ʬ��T�X	��@�dV�-���I5�b܊�+N(���y��[��#V2�����pX�/�)��p�A
$v�9k۽��Ш����I����D����a�������K����{i��!�}�`}�o��C�����҅��P���n����s�\n��r {�o͉�k�x�B�R��B�W�p^�Ư7,o�9��H�t�t�g��<�hv���4�gKMe��%}d�+\DB���l ������*��g��"���i���Y��,��X!���,	����C]��L���&�C!�!,�M��|4���᳙g+B���Gg����Q�v��[����kNNv`R�ON�<�L�
n�̥?���W�tПg����E�7ީ�0Wz��{�0��W"��uSi�[qxt+d<�gz�΀-�ku�.W�lf�zP�vLm>� X& XLz�?���^4��+IbDbV�ǐ��5�!������sc�(Tj�YJj���N]� ����T:9D��9$��ER�~�Wj�򭏀5�FO7�&�ͲH</�c��x���&�s6���
J:DŞ��1��n�ǒ�́0�6�1��oC>(���ê��u�K�#`ˎ @�0Ɩ�Ύ{�EM�=�Y˞�+ӯ���Z�.��X�UY���Z��A.�S�T5����.�j��aRk�����"�0���D�osڒ�Ӵ��x�/��IQJzki�@��_5�s�_W��A�z�b�D:�)QZ����m'8b��J��	l��:=�J�1	��W�cH�(Hf��Fv:t���ln�D�����d[�i�hs�g\oE!G��/N&'�����+����.��D��TՄm*�P��S1 ���q�9X��q�?c��Vt�����?����l��)`�;54@yn���B�8�Փ�W+�6�֢S|y����n����CL߼�C�0�`�ލ8�qp/ب��Q$}]�.�n�Ph$-w~����ƻ���C���4����?u���J���� �xp�%�y������0��"Q3�������'�J�A�tT����v!��OZ�I98V�Q�s�L�LV����>����G���x����a!�R���d.B4)�9F��IH���ު�I���#�˷|�����ia��k�|dlgwLSi.�|�to([D�ZKf����2	�� �U� ��c������ou�9ߔ�M�"׵�?"�`��蕯90�uP����� �=��k���1�e*\h�6��}:]p5��?�&�2�,�j��b\��e̡�C����8�Ր�|����!����։،�,?+�R��}}�b�VRP�D|��@;4����4ӏ_/eHC��E�VF��^I��7�C��:�h�-��/�.|>�z��ǹJ^�MZ����:��#�����	2�KB��v�������GN��P&��yQ�_���gȓ�00D>�ЂJ�����x�=I��c�׀�o�Cm���ժ��Fe0�̤(a:��um_:�����kTF�a��Yu�7<-Y�Z�hs�am}�#�����y2�[�=O*�*���9�b�Q�Y^q݄;f�����3t*g���ج��/��b���E�[4�����T�U5��f�0d����cA[mN����L�kW�T!pn~G��zXm�~
Ă�T�dt��ЛЉ����jy�ؖf�����CK���SXf\)J �DӉDHX��J޸H�	w�8�f���W���#4f���̆+�EuH�A�%HG� �K� �D����u<!��u�^X��R�B��~!њ|R��ֹ��bF�����QnP���˚�v��\]�3^S&���*��l�t�G��d���2��Xf&���G�?�'�߫�}Н�2����|���
���$�6�]�衙]�*Ąot��Ɋ%,GBI�V� )���x��X��h�����9=��W�t&#����g7=H!+V3��i�(�v�7;y��ek�������f0�]�P�p_�ǜ\oa��á��w��E�3Z�m�'D�Q���<ƞ��Y�i>�}�����N��Jӱ�_Ys�kK��~9��U���o����`+�>�P��'���Ԥ���˥�A��>���,L8$"*
gK���$cv������ƭ�pyr
�g���ua�&�G	ӻ��� ��bl`�9��_k��*�P�a�a;�ߚp����d
4 ^�K�F�� Q���o#�Z):?�����U��Lc���Zl��)NUer���F��P�pc.�tY����jN�nڭnM�-}�D�k8���-����^��XGN| ؠg���Xq[R'A>���)���(3B������Ӿ5�c�xX���Jrs �/\r� �������+�T��]�.���T����;U��e��u�{zV����+�ֆ�D%�B)#�HK�Ujm��㳈��IJg��Pӻ0f���E�2w��t χ�]dEHKؘm����m�e:<��������� 5���9T�}�Jjݘ�1#����~&[�#k�yY�Pb�~ �]*+죲���e��*X(\�ҴO0 ��S�	{G}�s���b|9KBbi��&��b��Z���h�Y@&_��a�݅��i{7[��z�(�h_�����|��U�@���u�My�nΐ�$gb�L�5�IO�Z/n�z����oS\��ɗ�T����Wm�z�%e�>A3������������;9*ޚ�b82��G6j��_�ݷ�� 9f����hW��yF����(wwO��T�m��ߠ1H�Ya$3��.į}ˊ��}\Pƽ��q�7@�FPNgOlݱR�(۵ݯp��8�
���p�� ���k�3�9?i��>O�1v�E��L�ۧj��V�f�1�g1P���	OlL��gQ୯��dY#�u���W�竅>GG�C���f@W$���a����~����2��������XN���֤�����) j�С���_�����/�`n[$N�L�DUY�gt���@�I<Nt����� [n��zbF��!,���&�!�܁�2I������;���Z(����nY��Rb��_�0(��Z�_|*y�a�ˬV����S���M� ��9�3��1o3!�K�����n�����b#��<���%�Shm�Ў�-`�s�0���cl���~t[B�f� 
u�wWou�6��*���RV�:��Ҹ�48����?5~sڙ�H�rE�g�|��U� n ~��]��xw����p��d��Sz�V���=��qdw����[eP������K��xo$u�ә��:�����qؒX���l��"bQ���;H�3�Ju5��H��x����IuŸ���DD����d�a��%���y��2dAd#\����Y���R���n@�P��0@�@�v�F�v8Yj��Zʌ����50l�n��|2t���e�h�eF��
9���ၠ� |,�VD��X�Y`��!I,a
v�ܪm��V���y;���i��Á�኱h[@�����z���/��F��Ͽr	F���1��=����މd���r��Ȇr���z�?~rQ���ַ�pP�����{�σc��b$�kȰ{7N9��:nĜ����$��< V��S�X?6q�p�.~�+����~�:��u� H~�c��:�S{+8�����x-��nL���iX^��ő!R�|r�g,!�Eu��~'���!���|���h���WX�!@�\R�i!�9�6$c()8� ��|�$�.�9s={n�UPG������?�G�k��1õ�6U.�/_���nc�N2�����3ԣ��4,'���x�[��fzA|��l8Ձ��y]964^Z	��ٶ�{��2e�`@���S)��Ά��fshHZ�m
�;���)%�+��!�(8��>�Tg��'�C��_?aZ,06_�d��Ѓ-сq�ȧyD���ʽ�țݶ^V!u�N����ZM�OK�T����{��[�ډ�:���TS_��O`�ߖy]O��%B@D��j��)\*����]y���$�|u��3��t�"9�S,�������i^�Y�Y��~J�.�S6�b�R�-x�1�<��>w�t�;�i�m��B�8�����P\�:����<W���E��"F���:X<%�iB�����KRp�zH����eY��]��#�g^��8d�j�*�:��C��`&ӥ�-+7@��$�Q�&Ҽ4�][o�c4l�u��{1�ȿ-�{h�aJ�Lr��l��X ��x������N6����-�Yћ�h	�D��ķ?�E"ZaG:tgwp]�H��d�Q�C�j�w`���u��}iDK�w��V���Tqf)�/)����̣�djT�S�i�����aC�I.��}��pf�g��舘ӉZy��֖�gz�O�k)���W�<�5d�iT�b���lo~;o �I(l (�C)x��F��CHk��ݢ�".dh;��^qy&�*��t�q�ږ���՟���UU��)�!}I������ע�TvH��V�?1��7�z�n���f�KD�5[���!,���#{J�8�bT-Y�碖���X�C�h�q?3n����X��əj͉���sf��鼝��L\B_�Y��Q��������:<m�s��D u��]���-q�0ko��&W_�c.
/H�Gk�k�>�H���&Qt?�~5�2Ui���{3#��A[Gb3�h����y馒��7��V.l�ᅥ|��Q�~c��?A�����-nZ��Xg�_��A,~y{�ɝ,%k*C��O�DO���]LN��_'�?�L��HR16�!���Ůf��o':.[t����O����ɼFD׫�F�Gk:�p�����؏!+�̅�1�E�uȵ��ߋ����K�����k�]|�4�<^��h�%�����^��$�9�4�r����d�5K�(Nݸ�P��׮QZ���y*{θ��&�Ԋ�~E�A���	V�3���9j���6:���g��eqq�+�U��'��,� ��g�]�wB�	Osf���{#�K�*,mK�d� �#�ǁ;3�����v_{�<���6/C'r-���{`XBw����F6u���O�9��ĩ(]=�Hm�D�֖R�L�W�D�+G�h���9�c�s>o��e�)dj�<)�x'�em�fd�*'`�/�!�L�E�l	�����
vN���x
�m�	f	7�j�'��3�e�z��֞�'_T���>��L�۠��������]�!�?���)Ӌ��zhB�!k�d��҅%hȰ���l5"bb�I�(�g�"IT�[O�?�2ɑ\�wD$E!�|�u<Ѷ+��f���8>)���c�Ȳ�x>�����d[�|dR�/[�vYy�1�c���"�Bx��pZ2�\�����:��8��+j�ޕh�3Y����8�W�v��Pz�iH7�V�GP�^��hMTSGG���K�:~�h߅ŢJ
)s��S�hbQ�m&T^u����Pq=I��1/�����Xo$W��I���q��EE�0B��{:�n���
�tc�y��"6W�C��xPG�
�FJ}8PYH�ĥ��ZRa�^"$���_������O��Ɯ;���1g1�M����9�|�;6O�ozص�O{��>�-Zr22w1[�e	�5Ĉxz�ќ
�'$�T�.����6����"F�)���ʿD�
���!��,�i1�N����=�,w��p�����R��.AB�/���|�oB�����q�y6��=Klx/������5P1"�����j�(]�%��s��E���9Ú�0��U�R�;�.AhZҙ�,$���u$GwD�=汅:X�N68҃��2�������%Q��g�c��' `	���`J	���h���m;L��;������W�&��J���w#JIJ_Hsp���0�8��'���-t�{�O�� ��7��S]W1W: 0�� ��}��L,�3p �p����<�����=��v4B <l�B�RCW����u�e� $sV���Io!n�!�g�#��y��2�2�6D�6/����A�� o�"�Z�w�� �m	�b��E�C�����P�$���|Lr�c�P�c����
�r���.�)�Ƭle�f�%d9D�鯷���@��h;�h�2�b_�/K���>(�.x\���Z*k^Y��~�!�A�E�Ѩ�k4�ľ�t��dOI��-,�:��v�|r��bQf8�!Y�^�g=�O��ύ� ���3�#1_��0�U�F���vIݐ�g���p��,R��k	�Ͳ���2���mn�8�>��ڬ��W�\w+�K+�����}2�7t2�3��
���[ze��j��.I~ Ю�5Kn�p<�ƒ�j���O������@΋-����q���R� �8O��ԴrU�X���d���$� ο�M����P0O{��)�,4c�0 �k%��)�V�������)DD��&����o�ݜ��74����x�䆾� z+��s~Ź/(�m�ft<o#�����g��Sh�j6x	hC���Sbj�o�,�X�����4ܖ�~$���T h-�sz+8��e=����Cg�6}u�O:�c��-��+Ҧ��+�[�Vu癛0E�K5�uA���E���ɑ�>�t�\�?.bځI�+y`�2��'��[�O�`qJ%���@��0�P��E�\q
���ԏ4�ŕ�g��yl�EUwp�秺Tq,�)|�A�nL-'�U�H_0~��q֋���@V�	4���ťG��͠i�(�ޯ{�t�����Uk�@ܳ��1Ʀz N��Ϗ�����kO����y�=\�_���cn�����mϿxİ�g�kF|;���N���{>c����L��$���YQM��n�1u�1t*�l�(m�ܑ�;3׉���l����y{(��\^���v���\U��Ǒ��ұ���k]Es�(*,􈖖^ m�qA)��2'�(�G,,tU�sI���<�r��o?�nV�����1h����i��������ib)%�*<�sD�.�փ=[�)�-#�<��b��)�!���o:鍄�ώ��
�6�? n�� ��`�[�ٷ��1����V��q����+�Ar�5F��Tq2!h�Ȳu�2����G4������0���{�pa�%}�&���<R�wϝN�
l��?r��w#{��jJSB%ϡf dya�4���ɶ�Q[�-��v�6%W^0]1�ݪ9,�Ҋ9N���;�����k��9��21�@y�g��?*�Y��c�H�m�2�Yy>w����ÓK��Ͷ|��7���\� ��C�P!a�3���8t�|-�bR�g�	� �A�͂�ʐ��{t�5h�$O6o� �N�����c,O[����g--Zp���B�B '2`�-�o�/e��E,j����Τ-.����f�O��k�W6~_�yR����r̀�H&��l,��h4���א���|w�(+�1�Α������$�M�?gJ�� �����z���Xd����p1�2��W����	I˲Q��~��	�)��#�W�������tHA/�_�9�) ���*/���i��Y0ű�B�F�ێp$�B�-Ը����4@�'x&^>;���;�43qv���|�V�R.-Z�[����m�`�b�>*���$�D�^��Ʋ 5V'�Z�9�weyvQ�`���q�PdXG(�b��1v�gf��&�>Y%�K�Vp�����J:��6�
��w��jm������F�d��@k�g!�c��=�x	I������,��d��^�ǚ6+�]:�~�r�
\�x���4�œEG�ؐ����b>'���K�Vb�>IK��
3�]
=b8��;;+���t�LL:��ה9q 
CWQ��r,J����r dS(�ط@/�W�K�mc0{<=��-$ۂP��*7�G�-���B�p`w),ֿ�褖�}�4OU2��O�ŴN�����1U�2��1�!��#7-/ l�w��~~֎�E5U{�\�A�h#��;����2�~�ө�ѓS�PwZ]0�?��ߟ_*@�G�ǰ�傀�9P�a%Ƙ��� R����z��Աyv�E��f���~yq<!�s�D4*�o֒��A���Y��/y��F�����i��o�|%�����N�Ζ~��-u�f�/����*p�6��X�B$�%6ƷV�7C�Bޖ!s�A���x�)����rֲ��E$���1�	����_��\v���s�o�?C� כ�tz0S�"��7��$':���e��T�L?y�V����l\�U��#q��BnF  �{�b�(N�WK�d(����#-<�>�.����40�;�L�$~:m�_v�/S)�7���z5�-��=\���R�9��i�8���������(�S�ts�9D�E-����	-����Ʒ���h����j�ѫzY�̢Z�\����7孂�+�~���6i�?��� �,xΘ׿������g��	rj���fx������g�"يG!�����K@��U��X�:>R�YG���癛_�`�.B�>��Ҵ��tKiXFR|�_T		�Z�$B����'��h¬!��
�j�M�7:�@5�9�,�����腽5{Zz���t>jMù�_Rl��ݨ���8��J�s݂��g������`�8ښQA�ܾ�OŀG�v4!v�|��:zJ�U(�a������O�}�D�O֧<ψ�/֓`U�S�9Y�����MpW�;OrX���.&`�	ŵ=�|�_���^�M3.���J�w����T��}z[1����Flm��D��%�y:� �=<]�W�<�l�	ZK.�>Uoy$��ԸɃU��s��������;�ۿě��`"IAgsiD�u`�~3�=�l�Vɽ"���t��U�x�@�:|�a�|�)�1ɖ��#�x��s����Se?�
��"0V�mp�t��y7,7%t3�(�mC�h[�Ѕ���Z�����11��>o��_��OA� ��0�?��.��V.?):[k}�JJ8P�!�t������fC�rj]�����AGS5�~�_n�׆䋲ʹJ,
��0,�nBfJ�tږ�����J�
��_���7(��݂�v���*��e��E�9s��K�Q�e�`�"m�VC�}e�ȬD	�5��#CH���댘J]+��^EEʩ\;.��SPc�D�M�.A����jmB�'�:��EIA;&p,B�.�ə�i\L>噀,�<�2�]�CA�5R�)�[��5a��������`�2�,R4#(Z�G�%�˪�I��������C7<��x�6�T�y5��r�3G�?n�`��Ϙ𷬰J���;��l��
�����C^��D��� ZE��h�;�Uͭ������F;�m����rM�]��]
vo0��w�z�e��3.�ю<BFJ�GP�K��[�N�+[�OKۧȜ�W$Y��Y	�Q~�'��Ѽe�(q����c!�&���_5�J�:�F��Nsd�<���o��D`OG�g�I���&;�ب��e��Ǩb�����t��P�����aQ�g���|�	�_ �~��+�����ߙ��f����-3	�~U���WD��g؉�d�rB�
X	� �h��8bw7�eo>ܕ|�Dյ{��%�ux��:����r��x���AD ��8�>�Q����Hx �.�.��(L;��G�yE��$��E��ls��=�/>��i��u�-�Ǥ������=էa<P��PآA�kL����YKe��3җ�	D�?^V����/�*����"��]���o쏡�����Oyy�R`͓ۅQ1�ܒٝ��r�]���Y��3��Aڒ���-?��S��^H{���SI�p}#h�����v�s`[��!NwDqxb��+�����8%s6�c��@'L��7��>�݂<��t����}�Ψ�&^ge]Nz_�I�rg,	�B&B0(d��E@{ �W����ȥ�GB�s����
�s^]}Ͽ�HA�������vZ,�Y\�cMAX���9��=<
�ȘFf�i�3n[�@ �$�ӗ���:+���S<��x(�%�w��!�.z��l�U�ky��YF9.�����K�}*�8�I���|dO��`�O���������e"���v`��w_H(�i���ޝ!��c���C�4�Ѝ(��?��.�"byG�KG5�	�؁��Y�����4d��sP����
ps�h�0�w��A�<���{GSQ���t��H6�9M�E2������d�g'G�[�!�J��ѱ��㎊�k�� �<E�_NrT�2���c����#���Ut�uE�p5���e�[{���z�܊�b���?�M�V�Z��s��H���,��6YӠ�O����
�Ig���ߑ��q$�D�P	��٘4���Q��U۔�����Ī�U	��Ƃ�^9�pP���o�Y,=s��T��Y����n�ă�d��֌E8��iV�!�0 ��T��ġ~F����k)L���H��L��Aʿ)���+Ū_W�O�Q�`�C@�]�2u�=��V���R������vV�	�pYڧu����JbT�'e��]_�JS|�$pwC�z9�t��A�Vgn�@y��ǺS����)���Ҙћ�����孪]�9����r+�_X��쯄�я�y�/Pg^	��K_��I̥��v����O�0��y� |'�R�6�`�UFy�2
3�q(�״�Ό�rÇ
i�Lc��(��w�M�jB��U�����,~l� D�R=;��rl�F�b�˥p�=��cֺ�L����M���;��1����Ju$FAz�����j����Bt~�)������JN�"C`��X~�Q2*}T�#`{GSƨ���v����R��
�f��݀�=6)�ԛ_����\�f�qK&bZ2��>O�\:7�V��V�'����_;QX��Ku���3ś
��������U�M��T_2����Y&�й��nT"�Ϲ�0��j��8u��9� wr�<����6���kJ���>��[X�b�Z��.�B���M�Vr��A��y�)-��7��;��4�=9C_��M��jпO���y�.3�Fv؍R��t�I(���(����T��L�����5���÷�)�K8�`b�Ď�s����z*D�]��1j�֣��P�S�[E��}<���q�i�r���D�ql2��R���|&�s��dx�z(] H�r�C���P�ҧPm<h��b��1����( ��8uK=��0,�=��Rb��VF]�,D��E�`Y��=��vu)p�l�ȵ}�<� ��u0C��?�q�`��#��_�i�%��q�W/>�pv\��k�}NB!W�"̽�Γ�!t��"��}� 4!l"��Lۡ�
<�����
K�ՌA$Q=,(�R�x���{�9�VBt�^�V.�x�B��i��w<H��{�\�Z �/Da5���8�d{�%��#�J�H���q�SS��D�"��R���aF�].,z���Wn6˲M��ܫ�;�d���UaD�3@G늳QgZ��z�,ebJʌ[q�{\�ֆ�U` �%j�m�Bݞ�LO��v,�!E�A3l�N�:R��Ar�w�Q i�Gd�{�g;qi�=4��(��/
�Z����ty�z���Pa�����z�ͲWI�t��4��T�Hzum%�!]3��دQEE���N�~so�m��;++qv��}��{�R���,6��{���(t틪�a5�Q	����ڨ���.��h{��>"�u���q�<�)k��&�G1_n�&��1�=ܥ ���P�wd���!i�Pa��r���%����'!\�;ܶE�Ѐvj2mfv��	[*��E1�JG�����	�!�noÈ-�H�Ĩa��>Br��$�m�������.�(,z��L�!�(�VO�<��Kb��05d�6�w���m$t�<&ѹr�xk����2� �a�H2��d3�4�7���"�2M�o�8�m]Csxx[_JGY��=��T2�P$����,yL��I��Ι��&}� ����m~� �
�خ����o�;�\��#Xc��9<��d�.�_�=�ڶB�RX�OS�(� Z��DGe�z�r����vu/��J�/I����{��k��3oƨ��Ʒv��F��B���]J#9K�P�0��Zm�Ҕ��oE�rQ*��J�j��в�K�� 5�����nG3t��w1,�^�e>`<q����
ȒЩ�$�4��t�	��ؗvp�������I���-�VK�Yw�Ro3	kܫ��Pܥ�\ QB�+�&���C��9��OTu��L�O�5���4y0O��!���2��Uml��pd{ƈah�?ܸ�@����j|x݃[)��5k�.1����hE�� �e}/A���В�?'�3
�x*�U�C��w�9�(��[� ���� (�=�ۉh�rg7�KT����fT,/����i����[s��]%e#�E|��ZH�}]:���o%a&)[�tY�3�̑O"��w�)y�����/Qh�6qW�X���E�|��Dng6)����M3�e+���:��t�]����=	� ��e����A\��M,��G��c�̄D��+��N�H�&f-kV�iJ������n�B�=�:r���tޠI��?��-�"�g��Z1K%	�覓هm�]C$�tW��(�ѵ�F.jJ�@��C�G-�+7iJǀZr!Vؾ|�󑤔�3%Ք�	���ha|����
�('k�Q�u������0$ �J蔡ۙB��j�syiL�7	����I[R�K܃X�Л�}��{���'��E8�
6t��oh�%"ȩ���e�&Wd(�`�^�3n�K����ܠW�(�l	���Yߺ����E�Ao:WM��2�/ګ�N��T���BߜmØ�RT����ԽT4���ۇ'%�J�3:�\HX�+�gzT�悫W�=kZMMY�;~c�'��bt���M�k����f���k�2�ZQ�����mR���k�OA6l�U��(k�*�v9���#��߫m�+����`v2Vy�aOSw1W�����6&e�;�[ %����:��k/��v��!��`�'9��Е"<��$���q�4巚?,4)D�����Fq�?��L�g��J	CV������b`p���[i��M�$��5NTs�B:y��|�Pj����8$+cc���v쾋�ܦ� �C$$}K��`bT��JH96���#�;���ӎ}�U�6����bKTM*s�|�A1}d;��q0zI��0d=�vȦ�v�.P���0$��?������r������v�>/-�ض��b��E9p��Ă���ͨ,<�T�
83:{�
RXQ+!�ʴ��@-�bU���i�'�~dJ�W�R-N���5�_p+��$��)�U�n�8�W�2> ��CΜ\_\:���}c~HfSӿ4�Zh�s3�ѐ�x(A���C�
���k6%yr��pm�@�	���TB��"�Z��C�_)��Κęi�qB7���{ _��)�,��w `=	�|�;?�ԟ$T���ۓ���d��D���AKZ��]e��`'ѵ;ɋ��#�o��{�$�"�*�\�P�hѸ6��B�]w�ϥ5M0��{�2�~�5���L��Q0����\tK_��d1-2���Y&��y=�42(mBO���]H�*|�����#�q����d��ء��:v;�J���y�l�V��� ew!�YK�\"
W���\�i�; �	�RӭPw"86�V;Op�c���:KlS�c��%�Χk���������r(FM�=d�K~�DJ��^"4�z헬��=5RR��)P���.	�P�S^���z­hU�W !���T����8�-*��Ė���r�[�;I8zF��pPA	)a�y�#�r�0� ��S7;WǠ݅5%~=b�#Tm�6����qe;�H���>�z덜��Ӹ�i�	:�D[�V7�̛=�"�Շ���-;��������Et�[w�=�L�Z(�Zj���S���e�=JۄkW^��n����s�橆92m𲀜I��%J��&��K���W���M�M	�_�Us����3l����=�'ƀ��"�bb��J���/D؅�;�r�a�<�� ����Y��;v+Ѿ*5��U��բGע}H�p$�S��� }�Jo�͜%W���:�*/�<|�P���n��|D�J-h}�/�$��p�(��t�� ��W�46x�1?����� j͵�1$��_�3e���eQ���B�ª��9���_��b�O�uܘ�(�	sD�c<)�BHfZ����bn���fc���r%��x��L��
�מ��\��������ѐA#�8�,�-��\0g��Th,�����܊fA���C�#ｌ�cT����P�~+g��,��+	:j L�vx�B�Q|�e�8��|>]^;0�359��G�~L�V���eOj��-���L7�0U�<���<�w4�Cv�CI��B�2�#4�����3j�T5m>M�|�Ȓ[��V�����w	>�>�����n.̸�����%��s���@��T�te�}����qr?�J(�'??��k��Z� z�$h��<ۡ)`CLjz�D��i"�����&��N��} Y2��;<��Z�pa��b�-f��
��E����*��8���Z�=<��}'���3�ǫ�[Nl�*&��x5���qi�'��s��h�>��8Eǟ;l̀&m�Z�H�͝Ut<"z%�����r�nH4��٤x���k�^H��G)&�����WU��H��)7���@�n_����?�m�x?*�q;�fD$�k�s�P�~��h�PP�
��p������ςX4�5C��� �k"�����Q\�[��9��sCT�Bh��c� C�����gQ�EB�8}�D78e���C*J���^�B�*"C�_+�ʅ�l0�Wؼ�S��KR	
��5*�V��[INdMu
��~����Bܾ/�>#����g�ā�
��픯�u�=}O��I-l�/8�+\�#d T�N�?L��2�^5�����=C�b+NB$8���c��� [M���ڒ�̉C0�����i�����X���L��hN��~����uO�?�]]��$GQ�'������\/�GIx�'��l�GF�|ojN�}J`�u��E e�爺��l��?`�_�H��J��Ho��"�d�O̿D�V�Ŗ1�?0��5O�z��p��G��\f�xv<<�2g"�clEWܮ�H��1$N3~V��`��cA7Db\�ɴ-u�2��h�t���(�Ed��S��t�wF�8�Km�t�Vtv�*6�a��S�z�C�A!�"��Mmu��az�>f�0��)g�����\�^^O��qJ�8
sV\�:O�*��y���k�S_��T�����!�Z������;����G�]�o*�S�xS�U��/!�_�L�v�ǙW�����]�)��1��Q�a6bCC�����b�5l��m�;�6����E I�}g���J�Lڃ�*�t�@��9�I��V�u�#è���q��:)5e��o�fOI}v��nu��B�IlB�B�1�s�N�i%ڨ�ݺA6��uL7�ݝ^��լė�r�k�^�P@cb������|4e�]x<LV������w�RU�����R�f�a_p�0��{��I)j�0C@f�b <��3���s*f�H������(ǵ.b-����ܒ"$;#�ݿ��;��z�����vu,��f�@$� {&��՘�W:̞9*fΥ�,Q��ީԐ�J<�X�G�{�Z	��(��ي/��h�?��N߈�8)�W�S���L2���B�6MЃx�D���W�#��tjI��� X�\��W囗A�ؐ��{����KlVʼT������.t���q�~=m�3k���(�?+��o�(^P��Od�~�Ji�4�=;]s���2��6��v��z�j"�P��П���EDU쒞��+�[-	aY�+#l�`�;�F��gR�}>��l��YNO�q�4+Z"g��u�#?�NA��4V��K��F^�� ��W�v��l��{�Ԅ�3o�����s���`�AP5�DIڳƘ�C)������|�ã��
˻JΟy2�_�8�f��K����'6u���`��*����gI�_Tdd����G������@a��[�K��L2�������}Hw��
�Mj(k��\0T��V=.�m6M5��NܿD��p�-l�.RZ�T�cC�����B�{��9%�q,e���N�âh�+���t�;Q})9��)]�c���
�-1�m��jPpy2b�gl�7�x9ǒ�i|e����.����
6��#�l嘭��*(�L^e�ቸ�V�6����g^����3�6���T�UN�6�Lbe���F�H�5�YF��gY���v+Y�P�"����y~j�ka3�o)oqW���w8zm�ė�+�=s�8�B��r<�cU9gH���t��ӄ��-�-yn7����9�a�_E./ʖ���/�eݧi���t섬ߤ�ƨ�р�I9���4�2�2��o|�]�B�d���5�s�*j2c�TyP4GT���tk��Z;hTO�ק���NCژ�e���>��O��o$_#��;\�	��,w��Vaq�-���s���N`�@dm�ެw��'�A�u�%�gєq(��G��X�v��9�l���K q�
�`m�/�[ְ������tn�� ŷx��ϊ��N�r�RJ��L/�HZU��!r�\�7!i]�d ����tԷ8�Gm�O�������g�4�.�[P8����]�������E	m�� t����Zϸ�O���/iٰ�|���"����օy���zz�:]�b��屧(��.��Pt�o��`A ��һ����Sv�r����x�}B�&o���&�d���������{Ŏ�,�X�����i����Mx��)�Ԙ3k���R)�����W���U�����u����C��U�*��hM��Z��E6�h��q��`�m9��.�i��ߒ3�y�ҝ}�Bɍ����a��W��I���M��'*�1����3����6Z�����`�.��B��b��7�}�5Ɋ5yȂ5������*�K��c�N։$�>�9�MO���f�����A�)I����)������;=D�PUZ5H��67�c3+ �|&M�1�R�0��ﳹ�Vx �b���0K�Zp|<7��2�'�g�|��۶!�A��'"�y��Ams�/��QW�%��H�Jf�¥�$���Yt5�%���A�q��B�x�Dd�T��t��BOƀ&8ȠX�kL�E�r��bƷ���{����?Z�-�s�XaMyH��20G�S��		�#1�w�	��*]F)RXL��w�k�Q���?�.\����oEisK��<�@r^�MQ"J�O�¿�:�
���;wr�0�̥;�t�J�PM�xJ�&���&Q�	�.ы���1���Ҕ�m�Ĉ?B$d
<4Rei����Q� ͋� �oh"��=����A�����d/�*�Mģ4�E����^������#]Ü������D�I��V� a�V�>�7���]�ԛ9,|�b�<�Q�s\H�Q���U�����*�~7_�e��9*�U�٭������m&*���c�݊��)�:��?�j���~|%���Y)yrI���4����ZC����4���bϑVe�|
m����'!���@oQ��^�fښ�t�6���n
��k�1��5��y�Q;"�K����.j4�ݎ-�ڷv]WT'���b���\ճ��\
/�i�l���8)�s7�
�vn��/h��"�< �P6n�S"� ��Y#�ƵD[r�!��K��� �0	�_;KߛG�ʘR�8��^d�V�	q��#W$M����#�lo��|R�^:񳎇��Ѣ��,��.�Y������N�9��b>�� )
��M��XU��E�s�u C9&�Z�o,���*}�?���*�YD4Т%K@�g��#H���qFcL�ch�\MeF��1�9j��Y�Ӗ]�a��1#�e���܏"}��88y	ǂ�<`\#QF�ڲ�i�:���h͡���ObT"zgi4~�#��ɷ���s��~O�N�}�چ��	��gh���_9��@�� �ZϨM��g����P"I(�_���_{k4���u�OrK�u7��O�-�s/[�K��h�$����f�QA�Q%��Aݧ9��*cY0��Uo�9u�͒�F���_(Ɲ���N�g*,���^��hz�.���݃[���4(�� �)B9���4+��1s��m�:�ݷxD���3�y�|ht�D�U�6-�mK�l�k?�~��6�~���t���mK��h��DH"	�Mo�b.%^�Hlz>¿c��'���8��r�bR�	pM=If�펟�/���e���#Eֽ䍆{�n)�<��B"z�
O7��)��<�5�ǵL�C<S�8�\/�A1}�Yl��-n(ΒJ�S��b)��>I���b!ԣ�w\�ý'N۽�V�dv
 5[�$�V����۱/\\�e{[#�P�������t�W���zo���٩H��������o*��^��r�/u��e������;�i[O�f������zY�+lN���"�%�H�@��\ �_� x�(�9��"I��tiA9i�+�*�'�������<�8�ęn��5--��Yfs������F��=�ܦvu�wG�T;,w(�1�jʣ:8qCt������g�zv�Ǳ*Rě��W���]t��x�i7-E��$��d�pr%���S:8�ic�@�>h�Y�n���i��zd ��\m������bݞ]�k��{R��5�U�$�
�����kLJy�7o�X��5`1%����?��g��{^p��b=L��'��ϻ'�4w�^9�~��oM�g�5�@�+��<϶�2�ȳ�(=��UX(�ee�ɔ�����Y��Ga�JC?0��-���&�Is
�bz�8�W�@5|�<�D��Yj�׃^V�)K�G�'���%y���b��G<w?��t�U�6��@�NŘC�1��D��fŦ5 \zKH�Z�Fx�a��`;'�L�ZQ�\���#_A��W��C�G�n^�Qу9>�H ����6{Z�T���`���y�q���D�L*P��_�
�tP�b.�!
��S�No[�&h�����2��7��� ��Q�	E�[z�ܟ�^�o���(~>��Ƥ�F˳���u�#�r��Ғ�t�%<XE�<�& t���X���`g>���/�(�����"V�M:��� �{�8k���W߂���qG:�%���2fi-�ʒM~��!�԰_:[�q��s�����u�PɅ�����
�3��}l� ��@@��_��!��˺33#�3F����v
ݚd .�</�h��ΠS�]��B:�l"1DZ��t#�J+B��}idr��w|Ȩٿ>��<�%E��X	w�N���>��k�4������7iPV-vs+�2�Ǟ���BW]�2�$�R<�p��Q���1�8Hc%���'�̮�n�[���3x�l�c�����KgV^��ͅ뮿�b�~���ؾ�'�#:(�^��z�?3�|��y��������D��˜C�!�Ĉ�~i� ���aT���c@d�sg�<�T͓�8%j��o���͟��\lq
^��3r$�� �+� YI�
l�T/���TxӢ͛2=���]!�Ɯ��2چ�@Q�>�+ݦO�k�q	�`�Ns}�7KM|v/���l-r��i�H
Wy�G����FX5u�.玀,�]kbD�S��C����0 0Z�$ע�ֽJ_�kِ��&���[h���AJ[���p+��D����=�g�ŰA�eE�4ys�ܗ�s!:�{t.�Lp��5�H(,��#��M�3hT��N�ǖs�B׊-���G�³��+*X��>O��y�w�!Z���x|���$#V8�_����ť���%�/�u��)�xC#VtB�`���8O���x�N�*$��"���nrO���C�#-w:b��X�	�C@�o��ma+a�
.,�����w��=gB�rD5����\l:��YL)>+k�_2.���Z.
�b�P?^�r�.�7��%���m��"EFm_WX���Me.��	c���}쾤�P��j՟`Բ�"�#�hNP��"*_!Z����=�K:���g� $'��C��"���F�3��/�03M�1�N���sc�fdx}1��z������o�n3'P����ϼ����8?�+���x��e�/,Z�SZ�S�j�#�¨4��?�6f�>���A[}ʶ$4�/��g�r���X~�1'�u�a�Q�prMv�؎`EJ�h�KZ[�i�d�J�,����V��{>Q�O�y��n<Qag��������� �q������\��l��>&/?qo�����4� ����6w�Ơ�M��F�����q�������`�6��v���Bؔ
��:gtq� �u~�E��ZON~ͳPw�U����ݺ�哦��:ٙ)@>�%�[�R����&$�Sc,�js�@�W�kU!!u
 2Z[sp��9`�zQ|�"j߳UUnV�*����4��㼩�(�=
{iИP���vm](!�30�D�'�����-C��2���3���{�j\���ϖ[���<d /V�@B��n;������Ⱦ�n�JQ��t/MաbP��y�}[0N�펀x)���J;"�.9�Yfv��3�A��H�H
���L��1f�.�a���W��K��j���CfĵQsE�����3��h����6�	��A����lRiw-KYm����7��	�}��k�N��5̄!���pQ��G!P��'\��9,��gވ���u�K{M���7�'����+	��K뻷���r�F�R�գ�P�X�UW��s�����@�95_u���m~��~�7���(v���߿kJl�?�r��<�<�J}8^��>ƞ� a֦�������J�~Z]�e��M���b�x�D����yQ�$q[��Ν��(�?�e��/>���{�-O맄6�`
�[f,��զ[f���jzV]e��h&Gt��>�b��mP)`�7X��3_�F��� o����QA�3Zb������v6vE�,=#e����.,�ݐ�k/ �.�˹��Kҥ}�����l!�rs�d�I�涽/�;�s!�s��2�T��'��R�����c�ӓ��S�᤮n���:2j��s�Q3h�<e:��Z�Jx��^��Ε�<�1fMeD�ZTK'g# Q )+Ĺ��i��-��!�2�#��
=��LA�iě�p@z�׽b�����G���Dk�n^�\<׻��2����e���F�?�w�-�#�륂oELwf!-�Q�c�K�7M�[:������x	�� �T� b ���N��!(��4PGw�ϯ~W�DxU썉�&zj�TW��Iy4�F�d���pW��YvF��e��$���^�'D�>�i�]X�8���Q�۹���y��;G�b�� 9̧��h�Yn������V��h#�nTc.�FT#�N��Me������5V�z&O��"�i#ϣe���x��.���ǟ��5����=�O$��J��X����y��3���!	����X��H-TO-��dݻ��?/����j�����SE�kCMx�o������~�,o��.⣋q+l
���k�S((d��U�OLد7�G�0$^�%H4�]�f�Qx*�)J��G���C�V*/_E��8���_�������)��Z ꬸ�،�����u�83�q!CTGŌ��BC��4��96V��|7��g��U�?3�<+%�f�0@��_N,�����X�D(���t>ʖ"�x�ϐރ�7��R[�l�BFC�i(�H��kMQv�@����Rz�i~�w�Y�_4�Ϋ���"b��ި�c����9��ȿG��աN�_�g��hs�������
o�}�\�Gq#L�=m�CQ�ʳ��ɝW	Y5=���<�X�K�'��M���r�BD�gMM ��\¼PY���Ne�!���?H���4�4��t.�i,
���VC�[�>�k>���Mx�Q����2�������<��6����[+�ۂ'�U8�ik��G�Q����E�GYl��0��tr�f��u9���K�$��������7=\����f��@\��7e��f�͝X�)�����q0��b �Y�B���sGc��Hh�bFS��	3���Bu�J����q�+�R���˙cv.D�(4���nЈI������T���s�<��G.u^���a��@���\��ɸ��f�F��|���Ɯk�|�.��۞�����l���1w6�X�~BQ2}93U?0ޅ��?�=XÌ�?!�kr�?��[Ca M��|�"w}����<[��D���YZ�IMoh��3�ìs$tJ7�fR-��ƌ�����B�*��.�7�ْ<�CM�J$+rs�O�b�#k*hJX����Fe�]W$[\I?Ɩ�~U����"�r�6�/���)N�a�q�j�D���SE��􀺞�;�u�䦩�a�Ff�D�WO�C�[��1uU.{�g�0������m�p��M<2�˻l����+�2��쨈H*���]4q~��r��� R�]����e���t��z�{�N>��sR˨�*TT�Z,Y���mw��?��"��M���!|�f_� |7�N�3e���I�z5���A��a�B��g��Xml��}�{\_B�O8Gj��;��F�����;� ��P��ybb����*���;K��N�D��[��e�|���I�Ң�Ij��S.�Ng��N�e.���&���9��E5�~��	��gYZO��B�k@���^ڜ�����\f�QD�ոp*k5��-��^�<����z�;;� �]�i�����G�r������u���W��"u����?V�լ���鳘��~0�N�w)���m����E�ŉo���{��n��on��8�J�A�)���uY�9֬��|t ��w�]=�f<cbW<��Kh��W���^[��[X�#��{��r���X�Y	�5�-��u�"l<��je�G\���=� |�����x��E�["A̗�z��ʹ��Xb��� 죠pq �@h[�A��8OX�G!��X�f�������£���dt�AhG0JH��4~���\���C �Ɲ�g<��t�2�E��E/���[�ɣ�q��r��ϗN�v,
�vd��"��0������W��!k�Ȑ���F�����'����Ջg�;Jl�v}c'�]��M"c_�>M��˾�����<��&3�V%��O����e��1K�O�)�ubj�ᕾ��>��ķ��m�W�mٍk ���5o,��ąC��K�^3\����QoE��?f���6OC��oU��Ʉ��Y��h2;�\x�R�k��[#z*x1Lt��&�Ō�2K2�!����^/!�u��>�JD����ko�"�;����$�r�/D2v2�%�7�K�g`˲�u��Y�j@SA׆L��*�ƹ�3X�?�*�����|��B_f�.=�o�����@����
��}�J�i2$�z�����I��̒B��HG��la���9����N����m� j�������}6��ğ��^�Y������/l�$��޾�Ў�|x|/éF� ��/|�?�ǛA��>��)�� 2��lfF��VߣS�����I�ǈ���E>F"^(�'��H��_�缈,�-571l��-Hޤ#�%��[���Qk�ْR2m�x%�Pfs�zܓ�L ���&��˫�xW�`*�6�b��a�k��V�\���9\��ac�j�=-/(�it��*�����$I|�ed.�a���[cFw�����yљ�Л[D8B$��dk���X`&(����w���+�~,��G�=�?��>��k��բ����EK�ŷj�$5N<�>�ݶ�z�8]qR�!�/6%��WiMB��7K(^�; �BTl.o�IH��a$�3F�DE�,nss`�O^ela�͍��0BJC���h���(�/o��o/Z�*���Z��>�����Ceg�j-���n�)��ѵ9VÏ�ӍS)�juZ�l&�re2����G0�<Bl�#>���%�0<���+?�"�*�����}]��Ի�@竌}�����8>�#m
��o�^2n�~�@�e;�>��;v39R�8��hm���'��'A��a�]��F��#�]�P�L����ᙗ*�L�{\-H��
1��+�o�V��FǄ}�I�KDl9<k+�Cn;�ђ�����=S���4�� �a@���f��\�vp���QF�v�S7�p�²�E;YAٝ�8�%Wck��y�ƂY�G��#����v�����L۾g�,�?��Oq~��	Ce~�ܜU��<�̻�h_��!�F��u���~�/���K76���x���,�R�9��yɎ�����,.���5j0ƙPH��O~v���<��Hb�azp�AV}�3#?}��L�<}�[ Xwyޙ�5�-=�3���kefҍTMPl�s	�%�ʝ�hsv��1���*"�ȵ�]�/��p��rD����LP'h�9��Qz����T����c������#Tݜ��(�a���1 Y�O:-�+��F�h� �勞���}~��eQT���aY�7��n��t��>i��b�(LζB�X�<%&�6-&{�D�"Zߙ�%2�-�Y0uGpITӭ?�W܋�~���$�D���ʒ�X�>��/�"+�(>�H�sj't�
�ٷ_!|���.�n�h���Vz��C�J"O��3�C7.K��;L�MJЏ�8��E)6�Ў��ꄮ.h
��/$s��l�i�DX?�i���L����K��6r�q����%�^��s�����G�C���n�f-��)����Ś�.7��(=��5�}!�W~%e�G���;r���=��)t9�41�Q~��/z�X�>�JhV�<=rST}}��-w� �!Gt�N�\i'S�kn�!������A�rstz�>y`h,�	Z�blU�xY'��^�A� fp�k�t��_��4��;��6�  r�Ҏ͕�Ky�����>9�UQ�>j}O��VT�+��� hô�*W�Z�)�^]�Y%���cIX�+�I��W��m�>U:��@��
//����W��A.%*�F^�O)l�/.�_C����DH��x~"�Dk2�{ϊ�)�4aVm���G7d@�~��+�k�W�P���>�$ �O���"6�繧>��Q��XW�~S>������N�~��~�}�ώxL��@8c�:c�z/.@�,���b���[����Dk1	r�l�K�Бꤻ]�띷�^r���3�Ǣj��V��y�@��u,Ԡߏ�E�d0�_W�K*h4���6hb �V`�����ż�G�x�U�_����Ϛ��z�+�����98� ��8'�|���'���A-� &F��s0��-�T����lStc[E<vG�7ՁL��y�h���ѓ��yj͡ݐV���F����/@�n���nk���̎���0��qFLK���,���7��wh�K��p �kx�'����%k +o�ͯd&��mh٠fZCC�Z���>F��*!�	J�%^�Zh��L[�N�þ���\�ps��J?.}͵܁cA�hg\�&T�Y?$솥��km�?��ݜ9�3L�>գfoj|R�#�%�)�Mո�v���^&����3����Z��$��om�lԲ�0� #���WlK�+A5Ö���~��2[i��J�R��Ub�-У?�T�����9n6�+�d�k�������7~SȻ�O���t�tm��:�C������� �v;����Y�y-�3�w�<\�L�?ta�1�7�~�k��	Db��_����<�R{��6"u��:%QE�IK��N)��ڝ��F������8�v�.{��H�YV�ѵ���\(.�	wpC%6��{/s�q���Mn!#Ǧr��U�T���5'3vax���em������eD%�%ʌ�"������hjr8*���eI�Ɠ��6��7��V���?��Fr��e�u��zd�2��$O�@��i<��t"��1��e���U�?��e9�a-ɪ0�h�\�I�'܆א;Ԫ�<x�jVTU�&.��z��7낏
INٗ����t�eK��h.bD:�"3(�w�_��&�{�M�.���������
&�vV����j�kG�6e
�]k��
;�U+=k6~�!�y��ܗL��|+��#�q!��_��a�VZ ����>ٟ�fmF�"����ޠ1��ht®!A�uL���O��(���x��#s@��x��,�ǽѼ��۸����� ���i�iv1XGeZ��0�xI+�i�9x,X�T�A=5�`O����Zδ���1l{�<�z.)2d}��I|p{F�����ށ���!S����zs��O[��C\u�4�ȃk����۴$�y�C�&p�P��M�ܚXt��+���Ě�E��7��
A���·�J��?3j)1���t߰�aTon`$��Z/G���$т��@�۞�6cZ)�{P�/w��b*����HL�(y����D����`�Y�N'���}����U�FKӡF�Z��}s scB�r�}�$E�1MDGf2�é�.X�q��w[\}x��Ӵ�[�i���m�P��'b
Ov���֟h+)	:tl�ϫ�������?���-��]s���X�/�ea��@�Hn�2�
�z&G�>�d���ʆ�IN`����܉TǩDbK_.-�_ 𶐭#��h2����*��O�A�?
��eb4��.ō��#j
�����~N����t��
y��r�Q��K:�x����Pt�@��ϗ����'����}1�b��
�w�$��1�6*T������Yu�>��0�����X�Q��� ��K��L��P.r_��4�ף�;�$!O���qTU���*�č���&_��r�#�CoT�%MG?le^V;I��Jb�t�ɽ��̧_� 1�
��S����Ҡք�,6�\����p&�4�L�O�\��)�U��5e�e�LM�E��+"GeT�n���[5š  ywm��)�>���?�ʟ�Gʘ?N�)��&��dү�:3F�b �#���*�,��>�s|����S}$�phB�o�k�W�Ⱥɛ�n#�w�����
n��M���=����������A{8�����N4�#�l��u�r���i݄���q$������^�E�'[.���Y�R��)/�t�C�̯��@t��6kX�'@(^2s��kӦ �!��	��aV}�'�:X������Z
��9��_����*�͠��q�ޑ���\U{�����q��nM~����a�̼s��E��5p�]�!�F�Y\�T'-��b�P!i�X�4���3����;�K6�Y'}��I�D�*D����ɒ���y�ǡ�]Y��k�Z�c�Ǣ�a�l�ܑ��X�XHm���Il��Z��	��v��� �a�Jv��;r�� �I�͋3n�tTxNu�m\m���~�D���f�U��JЦ{1:�s,Ge���5���M�ڨ���4fyB�w�S7�>�ɠlF4�|�� ���$aqv�FU��ɳݾ��RwZ��1����k�I/X�e ��U���9``���Ô^Ȯ��56��f�Gn�z����͘OL(����ل���B�<c�*E��(�~郹�����q���Z�7�&t���\�Y}�0��1P,�]V�{-S�����y�od��D�A��a�ɕ_a��LDa����ÆO�=݌�=����/�ʡ�@I��M'ܽ&]dz�=�t�P�ܤ��r��+��S	[��l�j)�\=���X`�iހa�Җ�
S�mV����(M;n!�P)�߶{���~)�&G�'�!7$;��O����w�R��D�뺹YQ5�
��4��j�<������f����hN��ӑ�3���Ö�rF�Q�^�%�b�d��u���2
�ͮ��W�	��4�ER���N�w\���:�T�� ��"O�\o�Y�Ip�� ����/�Im`|
��CS��蚁��~�t]�bb�o�@j��n�14+a�~��R3RZR������4|~�W]cS��{ώ�]�E���~��P�B/J$u9�/	|+��� ����|j��Q$/�n� ���!8��*�������%0�NY�F�ҿ{;�g����8�v�߷�C~D�L�?+�L4�4gHw �"��3A��T�8���h���]9t�|#��m[�@���U��|FP93q9��,�eH�&}-Z���������e[���:��f�Qd䊩�T�T�E���7��pʘ��O�\b�B�ڶ�n�5�%�|�Z�������P��#.�ω�_�~U�ȉ�F�Z`J��}�$t��M[�J�ʿ4ܠ�|`@�P�:��O�����Q����s���u��rS<�'�k=�+_���y�@t�p-Lr�!E�*8z��Yݲ)h(�,du�*�4=kk]��C���38b�\�A�KxͶ��:���P����J��c]�c/���ڧ�Kф�$�&_��w��rx^�����a�n�&
��eB/*2���n�K�����~P�EQ'��('qJY��_#�t��amne?c���d�އ�GШ"Z'��@�,�?a /mU�;�@������!��	o�A��(�E�UF<f��'|��Y����Q�,21b�i�ԞJS���c�3]�,(J��8�*"��֯ڮ�S�4�V�!�s�P��	ɧ�޿�d�Y	�vs�����΢�}���H��5d`B�-h�D�C� v/q��;\��Ƒ��װQ0'�m�ߗ���>4t��ۯ����_j��t��WٗrH���o�'a�x������X��s���߭�T{�( �+��ai������C�J�uӺ����Y*�%��Y 5}$>[#�0	1f:�P+ ��q5h�$a찥� E=��+yb	�Mr�c�y�Ò�?��)ek���nY?�r�co��P�ts��+=��l�Ò5t���Ǡ�z���*t�Ӌ��f|�{�������a4�b��Qj���Z�R�Bvؔy̚�;y-�'����7 h���J**�������.�JYF�F{��,��>�J���i�im�lv�;���cY��)A�菑���3���"yX��)}��mZ���4f�%�%G⬻�u|'|��|-��1�Mdo����D[�;����	݃�8V�Q���'ey=��=#�u�M�H8�,���+l/��I�Bm���d�I�q��@Cb�,����%�&�c��BљW�~��%q�p-�Q#����WEu��v3��Ta>���N��rI�{Ш4�5$�K7.wM�o��jr<�nJ�);v��Ս�b9�Ao�n���P���t_��-�L#b"��H�}��ʲtUT?>�l���s�3�6����-��0���������fD��~.��B!�J�$���̧��F��������cu>?�<�k&N9�C��G+D�8�WM�:ڒ	fC�bi�t+�"����⣄��/��[��Ĺ�Sgpw���[�=8��I�i'c1��!��ʪ�U��\xn1Z�#M�T!9 ^��l�����;`��pn��q�k��>ͩ���}������s �!�]u�N3!I�W
���۬�&��:`00r�����+�j��*�?f�et�j,w�����Q�%J$�'n-�͹���� -�j�a�^��m��6��2w��%D��u����r\ s;H��0_ˉ}�z���ܱ�����/G��=�U�K��ġߞ_��KY颀/�MF�ҫ����6��i6:G{�4j-�=������d���E�ʪ�@b(xA��ß�r�2�4N�]��^�Q?�&�,��lf~O ��'���V�qA����5�4(���xC�Wŋ��S+��I�E�/e����2F��\�0���/ �d#�7x�$f���7�eM4eDW꺱��K�P����E���ʱ��@Y�O&��*���l]�7s@m-��6���ߒ٧��"?Sf��a������c��S�H_��O�"�k�c��C��waZ�9���E:��J��d9�
j���5{RT�EnzTF�[k�*.k�%-[��Vg��g� ~U^g�7њV�8�h:�7�ߴ�ey�P���H	x�C��΁���E��?����[9���bNef�W�~�(D��o��<�;��p����A�Ɩ?R�����Nm��Ms�^`yQG���q��&Q�/������O�0b�o�����K\�����q���b(A׳0ٍyp������S���ɹm/�YaO[��J���?���U�\QW�F`[g�V�8Ƴ�W-���f�63�1�VB�S���f�����_��U�<,�jJc��6���2����t�g�2��F��_W�Z�ĉkb��?�)�ѳ�H����˸rP��B�La%5��̥UR��`�1P������G�<�'��iX��Ρ��I}�~EPX�?%�0��!���i���ہ�VDtJ.����,�2����To�*"���M:j#�����J]�.Iߎ�B܂֥�ǩKĴ<=o��m�쯻j��R�#�>�ၵ�ĜL۹/�����g_5J�H\��t��n�u��R"��,����g�dlp��y[3�d��Dg��>tV���e��	�1��3�A�N*�>���ZW�E�����6{�p�I��ы��S�w}�|�|��&����%��i&]N���q����dG�mُ䒒��o��4G��ٻ�P�ns��v�0uaMFԟ�!s%��,��>�衈��~�@M��T�2r���3��[]��rG�`�8N���0�ת�b��F�+]��@N�U`#k�?��K���L��>Dr�ʚ���D!	(CJ�3\���X��Xf�+w���`�����y\y��Q�_�xq�/�ìQ�|Y��0Aw����g�߸p���i!���_�R�4-�i{��hC�;R�sV��73au�u�0 g��F�2_����uH��}�gz��ÌA�R��NB=��$�ց|���J�p�U�E���[D�մ)���D�"��L�^~߽�r�<=Q�لB�A���������D�K-}��#�&��)&�:]?Y�%�"����!�;���N`|yԋ.֫��9SlAy�w� S�'� ������3��!6"<���y�MŊ�X����<�L�,�~�On諏G%�i����1.{4�{d�'��E�P'O	�R?�y�Lba��ߜsF��@�k���	]ӏ�)��u�.�ܪt�F�3��+��� !K�]]S����w���B��re�����`�q��Z5��{�%vF�}�P���5^�St��&V��ġ��,��/�*.b�i�Qz��
����Q:�s�IyŪ�@y�"N`1c<j�[���,�p6�Dm�����+�C2�Љ'{w�.���9�yn�wSK�C��	R/}�p��2~2>]4��]%SiNҶ��{�4�?)j�˻D�?m�z����V��H�r4����\�!���3n������k>6�����!�����W���)���:.a��C-0�v���/�Ej��� F�s��UP�O�j��2������RCd��91|+%6��&,�.|�C����0=^!H\y�ԍ�b}Q��P%m��u���7����d��� {��
W.8�3�)P���i�Ț���O��!v��tPj�K��r5��i�c[x� ˰�-ً���09�/�@]"iF�K�)F��3�0���|��#|�s� �袌���R���/�l�ζ3������1EʼMo����|��yOe�{^8��6�7� q��O�����sa<��vS�W\�]�=���5'򷆭�,�Ub�kjݻ9�sT��!�/��g����	n�;�����5s�9�_�`T�1Rh�axC?����T��ZY��#6"�|K��T��B�VA��ˣ�6&�*7�"�%#����M%KO�Q7IF{��[ta��L�B��y1hai�_m� �k��O�����ҿ��N`�:��C��<��������P�z�I�h
��7��i�kW���mwg�]��f�΀�$��*y�TP��w�%�r��#p��*\�Ę]A��ى�p�u�Q���v�X+�ٟ�	 "8Q�3���1�;^�^`Z!��h7�;��W�+�e��rt�d��1�h���� �FȌ�p&z�g���#}��`)F�Gfu�蒇����vE��"*i��6����}>�X��n���'nv�03"��i��3s�Ѻ��S?�S�w�o�g��� H�`������"�"�n�Ox��lц<de��%�k4tUK��=���e�b��}�o��Be*�'*W��lc��XA�?�a�d� ����d�Q���û�p�@3 ��dp�T���A�=f���@~0���r�z��[p�mu�ބ�S��L����o`aE6�E��ӌ��R�R�f.��	��:3م^�D�\T�!kz����4�y�L�})��C�'Cq������c~2�`Q=p^�=�#eiUT�����蹦��1�y����Mj�R�|>������X�BsĤŁm��j�d�����H�|�N�T�b�3�Mi��&�4�p{�n�?r�L_��/	h�Ġү�������Ǖc	� M ��i�\��֩5 �}ZAY�{��"z��`�VͶm���F_/B���'߫]�}Q�U�-�7�5�'(}���˱І!M��ʤs����LY��.�g�Mb�a�)����d�S[D=I?@�"����r���z	��J� �r:���I*�{y��/�2�?�I���ʈ�\��S
>�l_�6�wSB�^�:V̼V\o����}p��j�! �Μ�}a��4M���4��]�c��V���epQ�f'��Ao$參���4�$���/z��H0m�'�/6H� g��P�t�s�%<�!�eJ\j����l��g;Գ�/s	C�~�}f��\�4t��ؐ.[}8P�6k7vI$�����l����Xƿ#��=��4C�R?���³�D�5�H�[U�Ϭm�z����kg����iH��v��fLp�$T7Z��y_,0��2���%�ݜ��-ǳ�ǀVp�7��M Xd�?��60�6�yrz8�l����hٲW��������ZR,��y\�B��$H*?�Zld��B\%����-�1�`�+pGQ3ܲ1h/�J�^i�� R��p��IT+�T��;�p�v/���{Q��߱3�o��	Ӗ�����g�k��>��g��#���1Qy.���Y
��a0�����~����Ι�3�P.}��AcL�Ս���kP�7rjl|�?j�P�z��J�C��W�7�� LA��<�$uZ���,r].�~�7�k���<�j؞���k�%�(8^�!X;�VŴ>*�4�eA�/�L�לX*�3�H��1�J�9���Z䃗�h&�0�ݿLI�����M9�!��9�{����C�U���{��9���P�_6/�T����p�P��Xq���!-���٫���̨�32!s�h��NÝ-l�0��6�K�p�~4:ak��o�2��څǬ�ӿ|�.`����ڭ�cS�%@�߮1E���oy�4�p�{��	K���y]p�������y5�9`5:u\  H�G�Hy ���/�sT�P�nv"k+vb(�����(Q�� �Sg�,
⢮b��Y)8�`�A�&�8�������weyI�><��p����y�'���{c .�]%$ ���*�c��oQ$���p�r�$�]�}c�ha^��v����Ș&H���k6���u��r�k�Z���M<��"�2�'�"
�,g�w=�l��4�	sBa�=w��r f�fkO:�bx�������|�@�ӷ��I�8�J� k�Z��:\��η�v'���<y��;t�-�;Lh憵7H>n:<{�b�
�	��-��Qc�3Ǻ���GA��̎γ��6�"%8������3MY���� ��)��P{:!nM��?!�������P�cn�����x�M~aAV,v�q՝�U�lD��_ձFJ,���0-��!������Z���Q>�Ԕ>QK{P�6'h^�+<�MMY���Q4�w�X�LN~d[��4�zh�'����ʹ�,�ztV�y�;j)��ӆ���#��^o'��0�8�(%�N�,]n9��" �S�y6;S8�)��m>�c��>��y�?��� z;�E��~�.�� �0�d�ċ����e`gT�J�4�F ��Z�^D5U3�3/���;�?Z������L6g�$�R
˚j_���Iv�0,-�+�?���9��]�L!���x9cOY�v�&�F�ƃ���9��$��$OH��-�������u4��?��esacG�3�q��D���@Y~�eוR���eJٛ��XQm��Wea;i�ST~�mʄ�)�J�!�e4Ƞ"�s���Q�~�u��k�u�� ��n|���S7鐬�B�B%ͮ����	�m�L�h+$S:�#�,��vV��� ,e��ɀ�h*n���"��7�R��Џy����\�-�RFB}���Rw����H&���@���~�>	|c���s�_�^��Y�
���~��a0����8�;�q҇�C������3����U� y�;�O��-���]z��O�� �U�����o�Wjr-����8Qf�q|�JV��W�lU�"��F�w�*�a�?�2P�����r6����gb>1ŉ��.+I0pnr�	�O���?�s�8.;,?�0J��5_`���"��� ��^"<���.���l$,��J�,4�:��zld,$��a��̆P���䞈G�7/�J���^A�_{�Ɂ���w���y��^��G�:�����f�vkÝ����2���؁Ž��x�62�E���FdS
�G>�i��>��$!NPٓ���&��H#l�X{~t ��	��e�s�a��햲��d I���J��Nk^���lh*әV�Cz����6�!gAl�6C�B�9�r�li��"�b�V.��q���Ǡ>��;�_>S�kEx᫹�n���?AIY`�����yS�w؁h��$��2nXC�"����Z�l��g�ٷ��VgQ�f�� �B!A^-vq)���{;u�H�U8�������a)#J��������/1��Vy��ĭ��-$W��~{ٞ.� 6?^���q/ĤT4�0e���+R�2a�ĸPA24���l�<�봸b�3^�f�i ���-���"��S�f��v݀o�jc�F��E����&�3l�6ZNlSwj
������O'���=��X��&ā٫Ly�Cm��-���=��_�<�������ً���u��Q�#�t�����yg��l�L�`>+��FwW���;xش�������oa2kW$����m)�:ug6֐���pGzy�4�*	O]u�ߔ�S&v pu�Q0��M�
��aQ'���A�a]iQ�I���َ8r��aCk�{���v�c�Y?Z���R���u�a|
F�*�\�*췿�B�>' q���"ۀ��ؠ"ݯL��_*M��\��_TgU��1F�r�%�}�����o�L���V�Աh��U[�4	����7˷�$tzv�G���z�6�JX������' i�f4+~3?5�#A���_�aGV-�U2��b�Z����=/�j���9"���j)�$>�uJ��u#Y4砏1:b���~����g�IFf�̳�ڟ:3h�ϰߨ�-szҼ�=M�p��_��k,��6�7���"a
��?���;�f"�,[�g/BKh[.��D�����U�2Å
���?XI<o�<�z�E�ޟ�Mdx�S:�j����j5�P��m��z)��'5�p����~�����
6#�fÅK=Ķ��N]k
�wI4�x)�#�9�.5����x��x�0����¼�X�q��̉��߃�}Q��w�z� ����; �]��a<��/��$E��c���`Z����ԋBX3F��@U.29��{5=}���.(��!��n�Nۣq��m��
N'&5x��Ԅ`�;�q�\�%����eCU�����9Lm�jv2�X&V����N�_�[�H��z �Ʋ1,bv~.�k�*	�)A�Cc�26`��Zɧ�����'���E����.�o��)ुc�.�_a|��Vo�$%����/ad ����qEs�-P6�p1�z�便�[�`��v'�z�\����r��W�2$�OѾ�@I��T8TT|��6|eE�A�+jGMu͎�����E[��@�i�BuȰ�8��䝊�J �{������En�?߿n:�����tJ�Y(j�^1�#}nG����	O*�GJ�;�4��hA�U�1<��%�D-a��%��J���\z���G�%��I�.��oߟ��A��n�^J&�8ޝ>��Bz�p,���JU8�ܭhy��0x������t��S;������x��g�{m��!�GT��XOK��E��k[��:�B�z�	a�J�g��M��l��ec�8�vy��#�j���T��n��q�B��Z�vCI�O�Ӂ6@���'���L읋��&�9��ND�#���GP�Q����'�i�?��O��T�����3ї�d0�$e������W�"�|��S���dwr䝔�v�<�H���:&Sg�4߸�bR���~ĴV���%�̞������xX�.4ڳ���(X;#a�B}o2�}m�����H۫�*�����M0h��@�L��\�m�G"Y¬"`����?�&ű�A�f�-���f$�!P�?izm"��=<'�m�Ǝ�`�Ƈ�x�0����Ɲ����<p�q����J�3�3H�#b�7�$Q�^Æ?%� ���u_�|�:%|}\ИjA^�83$�S�}���5M{�#t���p =��O�&n{���0����3���tҐ ���p�༯t^������U;�f�+Ã'7��
N��dC���_�D���~����@��Y��i��Hk�)Wc�i6[Q��a����W�eq���f�4S�d>�8�r���@\�8�|}�g��7��!x������i��P�аU��R�����J�Z�@_��ױ�R$���h8^\��r�ʝ���gw@!�ΐ�T,?�l����e�M����81q���Gi.!���"��k�D��Ô�Ah��*p�B�?K*c�ƶ��Q\)��ì�n�y��y�J����fk�l*S�}&�W;���0��\9Q����ݢ\�qp���R��w_H��'~�~���D%���o/�;	��1,~�+�{tS���^�)2x���ϽJ.�3�0�zQ~�䥐M>C�X`v�=KI��i��s	K\[p�m:ŷ5~)4�9H�k���ɲQ������W7��r���9^���J��]� n�Y���<�r?bv��'�tW��<n������IF�p�f�õ���ķ�����J���B�b��2��j�N~.x%7B�Ĳ���/p|�}!���2d��ٵd8�J�����hŰ�����lR��I��ugxB�_EH����,���N�bX�w1פ��u�Ռ�o��>H(M�|��M2\� �
�q�	�$A'�n�'�#.��rX�|��َ{=��o�bJ=M��KD�(Y)~@.�Ԕ�j@�c`�Ԝt�)�����7^K�v!u���S2�u��g��[#;M9�X�� �Cq̙��[�W_}Bn�μ��?!1����MS�k��c�d�`�Q�r��o2�Պwrz�ݚU3'���������\� �tV�AaM'472�bg�cDr�WU2K�ޟ4���Sdrb��ꃁYf	��V��ks+Յ��*Py.��a��6�g+��z��������0O!í���|�\8���}Ax�u���M��ߡ��������Ns���+x[�tyϑ�]�a�����z!�+2|Ze���ۋ���$R�pF���/��M�I?��+>%����I].K�d
�,���Q�����4�䜱r�4@N�/�'�FA*�U����0N��go�-��0��]�|�������騹$}�?}��y ��Sv�8����-�oF�؎�6��5�ɒ"0��.�:��4,
�? 02�ܥM�$3Y���ڍU
M���Bveq�ϰ��c��cR`5S�@�b}S	ؔӹ9"4��[Ю�a�����{����N~�(�-������i��0���n��]�Rӈ��H��@_륺�k�Q�mJ�72��$�XI��`�l��p��cD��ЇEf$�c������	�i����aيѥض��.��\�	�ݝ�M����1�cr���,��J���������M1��5��Qe�J@�*�J���2J��Mx@'�NX���I��ˠ��QI�Ԑ�+���cBlf0�z@h�$���&��B�jr՜���$ih`�����N8�R�����#P]����7����pOt�	j��m!�xA&D!)�NK�'OE}�nF�w�9�y�(��?HXz�t��tT%1���>���v\'\�c6T���͚�O��q�kV��ZŅ���lM�!����(�6���[�5��ք�?�p��Q �:/`�N�����!,���v�p��x�O`��� [���E3�3�R�A��h���ī~j ��I4�����ξ�oV9m�^C��A�yr�Z��d,�e{>#�-g���j]ͮ^oF��
}�Ұ�5�a��x��*������U�6�_
B�V��x���$����<W�����8��Im.�y������F�{���*���]�&��&8�&�z"��Z����{�S7��E+����j��գ����|h�Z����e]��P�P��b���W��������r�S�穱��%h�W[��sms�?���p3��U/�L�^��;��)�����e��r �%B\�B���m�WK\��b�@}�-B��;�@���p�4L��'ޯ:�/��gB�	"Ǒ+��q�c��G��_�@�뇝���%�I�ȋ�f�z�~8��~����=��;UCa���9꾩�d���@')�S<$�H2!��eS	��t蔉֕��^��3��
i@�<+V����fk���o�D'�V��m����UL�ÖrW��ѧ7yː�E��R���s��c(^,:���(�Wwj-�/E<�"��|�w.�8��|��f�6��>&��LBxl��`	n+�VLJ*@�pq�o-�a�J�Oq��{�~X�3��j�:X�Y��'2��R4�S�Q3(�y4�n��)��sBJ���knU�q�����N����qX�~P$A�������[ `i͝�,�P�WҏM8K�5�!':M7�;^>��w���	k��.�Z���6�5�������O���>��-��d��#(M�_�|N>���M��z��=��	A*�Ͻ�D��V�Oz�����	ja.G�2�H��1�ݒ�C|DJE�|=���G�@�/�PϘ�
����P���a�.E���a�2t���Z��� �Vk��뭷���:�-��ʤ�%�h�s�����S�,�r��	2��O�j�߀a[X5�ɂ#��c\*��:l;a @
{^fG1�b}d�x��߄��֡�c��[]��tP�������$'|��<�d ����y��Š���Az1e��Qs[�d��{����LEE�˧�'�bc��w=�z�&�b�^�ʘZz��u�|]�/����c&��N�� �[G�@���*�D���$@�V1|�=	@�S�5�GD�#���%��i�zI���e�K��ؒ	o�Sxx�JY~��/�o�I<�=��8� 8�(=*�;e(єa���6ีw���s׹�o��i�l�G��Oa=VV��щn�����p��5o���$v��iA��V`9\+_t��é�z��>�Rcz�n��\]$�����fp�a�ia*N��}�`0'$tgr����"
 �w����eX!��p��M�W:���䦋��^�����*��ݴ�W`^�L%���e��7��$�ie�8;!'�����é�ٽ6�걏I�Em��I]#��0�����W��S��b]kn�0,�L_PC��4��E�Kh��-[��t�87���f(ԫ�������CEX\��i-h�м�\P���	M�Fdk|C��X{�1�B"�m��Ҁq'��+{C��R�}�Q/_�W)��m��ʳDA6O���N���A�5F� �T���*=���L�^v���Z��&L:$���.��tF�4�םIȗ���N r�N�J!?��J�U�N����sj�ԡ*a+D�*�-�č�	�{s�B��l�����ab�w�C�U�/�q�
X;�e'�O��|��vߐ��c�	�U���CP��ѫg��%�Rx�+.Xm�x%�b�#�rmpBt!#�p'�=Bw�2��:|�J���^���{��Lal1�­v���?��1'K��"U��j�F�������Ы�j4���Ux�c������U��l����r��[�6�#j���Ef/����e����r��+\Y+p�
h��=���芶�BL�&�u�({燔���ݮY�f�Bjx
���T��F}-�J�M����+^sQ��K_�M5~\����	�J4���Zsg�.���[	��W���פLSc�.�����QlOۏ�{�	\����;������)�5����X�W�t�V����r����O�-��2Q� uh�qrMuk�qzNQ�����X��qi�rs�3v.^���k��#��>7:*��k%:O�Eb�~"��Pe7���H��=3�n��I;�fՉ� ۰rp~P�����oY���牺7��~g��,�=a��L�M�ʳ�|���w�����叿�����,6:���E^�YO��Y
����#(	�s�l�N����v��q�}�䕂�Y�"Y����k��v!ջ��*��z,�5.���{l����!���Nf�-�r}�FL����s������,�}�����@���i���b�hB����i���I�8w�H/(}+[��v��őy���U.�@�K-��X8�s�al��#��9�(xb��\��9Xnl���|jq|�^�������:��M<���%���'��5e6�>���^�;%�ʵ�'�EL DM��w�ӡ�K�ֹ��RxW�!Up��5�%rI�p�!G��'���T1���y�V��d�9{e��9e��I�*~�h�X��J����<s�F�o�/�&p��I�x�kyQI5Jj�Mj���F���Sg\R���y{��u����y��=H)�T�$b���_��]3@-�����s�F(��S���3����G����s1vu	yl�,�$�;��l!G_̈q����XL�)Xp�G�X4mX3���8�*�����H�w,����eps�h���� ��#�) s���M|�`�ݐz�V6vǥ��|�/1�B��B����;�;��1>���7ً�y�Ϣ	]�8x�uu#�G��:"BB���^�}o�oG_���G��Ov
tZ�B ��&������W~U��Hʻ*V�%�-��W��.M�-����z>72�S��X�	��y�c�	uE�CJ=�v2=���t�B���c����*v�c	�u������F����<:���0X`�C,�b������C��B2+��Zdă���^��}��\q4�^{�A&����)�s��C�h�J�DO�#E澖zWdf�����עR����ݸ<�c۔#wN�����3[�E
�O�,� ������
A������V���A��<��n[̟ʮf�� �D:La����gSbyT�e)�=�������V�6(�M��u���N��*��b13���pȴ	�x�.;�)�1�B �kg��Ð��1��H4?�֘�?{R������>IzX�G�$���K��j�^���ZH /%���t���jj~��8��I�98�	���Z(�8�<�8�\	2M�v��<��󏙦����$�B�!�pX�Iv�nQ|�#b�3`��wÙ��G��+��:%�u��J�x3�B�^�{���"��P~t>,��(�;*`����#�.eJ�½��=a�҈B[���F-�cJ��"���*�������WzBdK[�rದe)��i�����.�  PM㱖-���&�1#��M�㳲X,6������S�I$�,�b���L��0�Q6`����*�i]62��V�A�N~�]lF>_6w�p3_��|��y*#ߡ�,�)��*1�#��^��5��R��k���Q��{�"�V/�h�z�A 8C�V�f�='�zr6՞O���
�鈉4c����� v�v�V���GV�G0��bf�kP���iw����hC�M��0�Q�$�;�i'�"~��S��шoɕ���"Z�]>��=$���-�h궘�6>=X�M������Ҥ�c<�_e�Q8����2��w�D��Vq��6������7��E	#�Nd�	���P�R#��DC����Q3I%��~�މ�{Oh���pI����J��NH瀻5ٛ�ìڤ��i��y�+����3��GK;��<gl>2�Q�GĆD�~�(^�����1�+�s%u��픧q�E�	JRj��լR�h�@|}E�q�Q���6�J��]]�P����/ŻIx��'ⱏ�&8���M)����X4=t��PY!�O���a��0�/��U2t�e��hgNH�6Ih��MhCR���]��.�]v�����g�Q~��;w�p}�����$�%HM	a�e�F-S�,%�S��4�T@8��<{;���d/P�ʞ#�!��߳��!�]ڧ>��$O6Ѿ˳ol��Z���gU�Asj������=1uC��xyꙈR3�t/l4`p91�z各���N���Sr�	/7ٴ�	�^E�ie�Ҡ�Ͱl������gw�V�sk��p��ou��2�,$T�.l�9��d���y�B����L��5@��X_�^��L��n/��J�`r+:hs��TR&&�YӚ�.��)����]��:�Y�b*�b��ݬ��`yM���k��@�k�yc�7+�T��+�6�#?�A"%�1gE[z��OTݖn��GЖ�42�����L�&��/W_�yZ�������P^�hM�9.�;��4;�i��zX��M���޴[��M�� ���{Q2�5s�N��lb9o�0.Q|W!����͍#��I�!��(��M[�?�s��ޗ��y�ku:�'yuH��8�-1~�(�����o�
���ϧ.�rP�M����q`mϿ�O�y:!n��y�	EU���=�f��� `I�%�#����D���-��2����=��߉Ȟ�Fnp��U1����D�_�~O2���%F~�Z��j������/�7�^�G�x�9�fهJ�x����Y�)1�{}A���vr��8�]�Ѳ6�BF0)���I��f���un�Pn��w�E��w���85����`.7AՊ�,�'�)8����n�ŋiNI���j�Ő�.�l�'&��&�h�t�'�y�#��	�1��H+KN��=8�\���c�m4�V���R�=��U�{7�*�:��<>7��E,�E�I����fh��EY۰6����N�$0�뒻��I��Ó#y�ct�R��7^����<�8(�]e��>�@���z˫:��v�zĪYn{��� ��YQ@'d	��=U_��I)���B5^eG�x�����m�|S�	?�E����^���e�ߡ�R �!n4����c�eT�9�,Ѕ�є�J4{PͰR���kJ��"��;��b�!`�=7(=��&��[6�,	��3|W�O��5t6%��U��>z:�#�k��fWI7W�qL�!tVh�zɍ�O�����{�R&�y\z�1�����t���S��C,ș=U�n�
�V*z�Lq�la��y�y��$��b��Y�Ͼ���D]��� �F���X������ӹ��ȧ�+����d*��s/C�E�3�����Ķ�"[��e����l���q���}�v<"�n9}h	�-���akL��z����~��m�$WW�*镎��B?�է/zF��:�i����	�O�]Ug���4��,�|�]�d~��Ԭ1g�TMv�����g��s()A�X�T���5V�2<f��Fb)��O�o�*t�}��)��mU�EN�m���|ݪ�@ƴ���87P��| C��y�Nl�^�^�ej��9/zE�� ��6��"�CV5�+��*n�D���K:1�������?y�s6�X�/�(Fs������[3r@R-+�V��G�6��`.޳������l�g(X�����~U���f��Y��X�s���*l���޹�OH	������-\ U��(�@@�I���V�}5Z�/C��T�����i�d$c���C`)y��b����t�������6e��y��x5򣮶�O"at���ȓ�K�j#|1�vr�A���	���b��-WM;w�����IA�Q��4	�1�榻����ԧ_���t�ڣ��/N�[-�鬝�� ��'���ְ�Q?~.�[p_5x��}��Y�r`G�:�2�xP�3ap6����l���9e�#Q��ƔȮ���i��-������ޡK��a��֯nl)��7�R�	e3��VjU`��7�YQ��w:۬1��"�艢�_a��̢>!�B�{TD�Z5C����f%QXۑbwB�Y��Ue���M2k"� bM����.�1~��R���� #�֠`DV�;��=�.��!~h�&��yvշ,V�'�� ��*��{t���&�Z��p�&��BRH�۸�&ϝ�F����BC�0�����6���4�8�$b �a���i[إDp��-��r�����yb����p�=!�K"�}{SZ�c[:F��f����ܻ�p0
�g�aX��7W8�m{3kU�wd��TO�D�V=��7,:�x��T(��p�mzGe%�kL�h'P�A�lAG���Vc�d��z���6̲�ש�$u����/��
:H��?x�����w�=��\E�f���R���>�(��o�2"y�!�Y�~HfͻD�Y�D�0��x:X`*L\~���6�2 ���Se~]��v�,�r{o��������^�bd�p�1¾�,Iy��:�U0��]���X� ��_
o�Vr�[���w:����O8m8�q��nlE0��%��� �w��l����(��W�d��q�%����/3q3C2�ڱ�����*��;�m���<-+AUI#�^ٓ�1ua#��7"s��&�M����\�W{�vG�P����U�0dL8k�_�Y)i��p�+�)��W��|ؒE/��`�9~�nx�𭟽'�����I�{,$QGڭc��� ���:%�~�ףZa��Z�Fz��rS�ƪ��	Q0I��t8��M���ҵ\Ha��E`�p����r�ڬ��n3r�_�U�T����VIL�yOg�|K�F��������E汞)�M&�?8���4 *J�R�b����DYO��W��R1�.=R7��Z��D��U��"�\/��̮�4���̌긔o|�K�>C��%j>%D@��U����P��<�^9!�b2���XC��h��^AP���\����$�`~�_I�'�O�\|�s��A��ڶݩ3��cq�4O���t� �s���З��k��8q������z�S����kP�n�c�XXy*�9>O�Z�Y,)CP J%rL^�	��`�3ڠ��!��us������*j �	��dI��N��Y�R�f��ڞ�CYZ7��-���5��iݺ��[��j�y;������UL0��>Y�o��n�^���i3���.I���%�\�!�MX�i~+{r�'虦&x��.�J��,�hr/�1�dK�b "<�n��bx�Q?�'���*���\y**�YG�10����q���*�h���QU���r�ͯ��|������W`=t?������{
���,�M�=���:��}9��w^��Q@<r���G�s�S��Ho��A���$:#2�I�w:����+��)	@hfFa�� �Z7���}��}+��0�f������]�Ќ�������55Rۑ4yU@��qu��t�骵�r&��6>$��B��,{�SD��:'��B%�#��������/sL���>'��Z�y�[jz��\���/�����a/��	,S{�M�_��]3 ,��4z�:��δ�Z���2q�:3�_���Ni'����V�Fk���I3�j��B3ejjphZR��}���d�u�cT����D��L���80%�HUC�=Ig��S�NJp��n�)�������WҴg�.{Iۤ����K@�^�h �a�J>��!d�V0�:POg_ո���Wn��;�9�|�̬���	IJ`�f� .q:��Km6D샔gTDE1d^8y�����I����6�,��%�!��C8����*����҆;��U�� %�'$6����F�j�3��}�'��wI�&���!.���`c'��v~�1�܍�VW�o�GNV�=;��yS�1�@�f� ���R~���u�6� Z�!��|��Ͼ�UV��!�@���Qh�{{��t^��7��	��k%o���DI�H�Rx0I�h�s1	u���(O��C]��Ҏ5ˆZ����z;q�����S� �\�Y=I��S��$�t�W$��H���Fo��qGB��"W�����iW旼PYB�;C�S�}�J$��~���r��f�V6����e�E�z?.�(�(�e�-x�h��ܲ���d]��_xι]��ٲ6"�$�wb�ܠX1U�k��r a��r��m�P��v]:����NOhG�Q&��&���㑫�%�������Vy%�e ����?��~�R��(�=P�#�;�[ ���D�~E�m[��Px�犙!���E؉G{.A���z=*�6�"�&��jH/) �]��1��!ߙd�����$��r�"�Za�Wf�}��y�Y-�_Q�ngz[v��g�֒yW�����gR��z �|�p�U�X:0.ى����^�d��$��o;�٦B
�Ͱ>|C�+��p+F ׼"��{�U��W�o�p�ž�%������Kt��U�Ѝ�o��UI���@[M�)��PU�ȉ����}^K�k�P~ϥ��^ۖ���sb�9�WЮ��#ӭ�be�%��Q�$���D�]�Ø�"�\�rbW�(�J6*o�y�y<vX�m�ɹ����i�8�"�y�]X=ۇ�<��6^���<����:�<�9=�E�z�a��]�ڤ�m�8ڼν"�gÄ$����̵�B��[����T�@������v�� ��a��$�6K����%q`�&`��D/�0�%\�~�^��y��>������sשvi���~��b���|�݈��6p�A�Kr;9̪��]���YNIC��Rv����ʙ�'0�o�n�L���H�׋0�HVh�Vы�x�-�"�29,q��(�k��ۋ�.�љT���2�Ө���_��ǣ|a���\�~I����ս^p[k�5�w�_�'ٖX^1��A�i�^"�32�T���Y��&�Ŧh�'dr���Z? �.ƛ�n8T���M	-0k�to׿ud�(�n�lD�ȣ��e̓/	�-�kL���qm�(�YU���ަ0Y?��>�9�E�M�A�"|�u��J������
�A����\0z(�fV+�L<�@\����o�������O�����n�/6��p<m筑��y@4�����aBH�.,z��i��Q\6�X�s�jN��'���hEBմ˶����p�@�3�:fNZl=��i��P��F �x���v�V	�w��RW?�����u�"��~�6ZAq�1ma���ꋢ��hq8�{��X�ׂ�+�&ߡ_��lj5GHJ6��?����7�^�:_т����PE~tx��n'�I�����b�N`3C���k�Rg<A�\x#�s��,�c?�2$1U�F��jm��kOO�~O���V��}�q���	8T5 ���u�<��t4�i�����'|~b�݉i˛]@�5����)G[��C:�ȰF��Dў�Hr�J�|��t���[2[�W&�K���ʛ&���������5��R��G+7��Z�B�� :�l�)�p��f�h5��ѧ�Qmk)��k0:a����C��*Fef	��M&�0�/`�J2����wڣ��L�Qh�1q�e]�����[_c*��$гfcKM��7��[P1�^���l�z�Y����qh����B'S=�5N��dO��'���O#Y�5庤N�$v�m1�ʃC@�]�x'~؏/���V�Q�K������0�V� EtB�}��B�$��M�����K즓	C�G9�6����y\T	�[a	��M_ly&+�|����	w��9�)|��+q�)��.��m߷��h��9PC�@�Nx��y�X���]d^�������ֹ��e�N�}aq;;���;�&��|
�ƾ�2z���u[���	e��m�d�dȉO��ts�;SV�P��[���~i��b沱��v^37�P`7Sq���еDg�t��m��B�I&�C�f��/[��z6�</���t����ֿ������m�2�im�+(i�Rv����d_9�G:9K��"������	75
�,��S\r�3λC��~���^>D�4ՆY�>4ñm����T����0�Q�M[���/&H��%�.�4�UJ���0��q���l۬`?��QW��xp��H����ʵܸ��I����F�rD�oE'9݊�R�&�v�P����McG���X
��l�5�ĕ:��Q��x��u�/Q����O�U��lA�2E�����a?号�7��MO��/ ��C��:qmQ��'��hڞ�`�#o3)�qev]���80UE���/�29��Z�`��W	9�W9�;��Z�Z79��E}y�OD�*#����)b�>"Dҡ���Y�i	�	�r ��yNo-<�hbp�5�bz	/#��/��
��Ҳ�*ӡj���6G�ן|X'����C�V?�В|�N�J�]/TT�%��>H�.�=������a�$��i��NҐhFݎ�ߵ�W���Jh/��'�ek���{�&�M|�
�]N��:�����g�m�̲4 i��̯~evX�F7� ���y��R+T��]��n�����C���
�3}�!z6��-�E��>��h(B$Ζ[�9�F���]Xb�E��$a8�hi��[�4C~.E�#����9ސG�@�5zagK����U�+zo�iO�.x>�ࡇdb��>����h�}�� My�.���*�Ld�跠�!(,���7O!O�	z�̮�f���eni�e]3di���,,_�8o�%U4'��9˘�|��ln:r�)���\C
�/9[+�S
�K��:�N��`{�r�c�j�4k���h����3WP��_S��|
u�4r��c����l)��mӦ -���4��I����B=��%��G'$@`\�(=Hߦ�����HQ���ٹ^e؍Hמ@�k��xF��?���cC���{{�O A.I�������z+3��KV
�2n����`�;�J�?�v{gH��f#6�I�4����ӱ������A�a����L�Q�*�r)Q-�m��E�?;�G$�����3������'b� 䩗R0n�ϑ��!)/<�� �F�nX��mY�
j�X��¨y�Ƥ���A�
�B
����Ͱ���^�4�a���Z���-����;=�������V,��ӊ����c��LJq/��Q!��uy*zobt}��>8n����a}f-c�:E{�~����a"'�w�hN�_����������N�?�;wȓ�Wn�'�m�L�Yd��&�/C�,��(��.>�h����@uΦ�*��x,Wz��LW� ,��uD�@���x��1}/��[be�D��R�;B���R s�3ݴ�Z䀌���*x�]� ��D:͆�Ra'��L�Ӗ*�Z��G�T+��`�%B0M�}N�2d�b�\��_$���2�E�[�\2<�v�N����V�?0x�5�oN/<���f�H�A�@G)��'F�se�[gk��xTD�+	���I����e#W�y#X�e4is6_ax��ͽ��S�UṡpA�Z�<O{�s�Z��`g���`�ɲy[�p��M��cK��%Vt'��+�̲QZ�B��D��Q�dt�Z@�9�_A%pd�,�C>[�8�:����/�<ŔpAO&"���pg4������>�	rSA�8x���Z%���[��Z����2���Rڀ�4�Ѱ-U�	�UK�Yز�Sg��q;X�9<
ٰ�AڬӘrZ���Y���ANn�.�ON���a����-�ʳ��?nUSN	|�;��b�F����?�Dj �vO�1��C�\s��4����7�֊>m�ٯ�:V4�g��F�l���;�t�>!�<8K<t�Qܯ����+��LT�4
��,���R��º=3��uJgӥ��<��d�Dd��z< ��!:D/�c�\|
*�+k�A+,O���B=�Y�w�i$} ��k_���F$t��,��7]��)���d�o�
��
�Y[/�������gK��֫ךmƺ#+=��ۜ���R�L���<�UW�A�(�����89���R�n%�B�(�=t��-"�m�Zw5�oK�;���ft{�ȑ����ӏS�.?�}�Cwh(\H<�UHD�k��k��T#��P{��^O?w�B�x��q�}���K;�%��~�Qw�4���B@�u�g^e�����H �����3���;�û��]��䫡l��/�&|+<@�������rW�g�X�n~�Nn��ɞ&��s35C��ƅ�GE�jdd(�m�����co_�k�t���������/O:�U�QM-2E�m�(����8*�AS5���Z We�/?���y����gM;Kow Ձ�-�������?��S���{���m�X�Wz�k.3��X��YЛꊋ�G
��|*ћ�"�T%f?*P-�۾,���=L�#����pG�al�lo:�R%�"����0 �^|�g$�"�4[2��Q�{]x���o�y�O��1�9I�����?YZ�WMzڈ���
e� $|���N�{�����T\����S�sX����ˢ�s�os+�cJ���
�1���K�b�b��ё��d}B0��(�W���-�Abe[ Uz�AY~C�X�'|��Y��"�e�᱉���yhV�ۥ���-i�oD�U��e&��&��Ѵ��D��bkl�Ҿr6:�&|��;01���b1O瓩i����#�DgP��(bL��8�/ED�𹄀C_,�8�Z��ĶY,�XaG�W"ʫEl����&�H�#d�%��]�:{6�$[��os�8c<��Ƕ:��f���}��=��i�E;��k֒���n/�g�<KK+��Hh@N�%��0��d��m�>Cp�F�o%-�%%���Ý]n�/�vЭ4��D��E
2����j����h�y�n��v��O�톢��@.��3~XQAC��K����\g3�c]
e%^�ۘ=���L���4 }���$�����AU���F���YS�z��7V;;�%8��m�~#,ț�rh�d[
e�(��ť�s���*���4�2��E������[��"���ħ��}���3�$q��5��u҄�����?��f��Q.�����$�Z����DI3���������/����Y�Yu��o,:�hSPԶ�2Tm+�X Z���T�7e�G ��Ȕ��m!|�X�ʺ3m��V&�F�h��R%�{O��D��ɐ�o�K@7ڮZ}�r�|�kWc,l̤ƙM,�O!�й$�Vb�������"''�o�*��Q��Q��id\�}=�>�L#@`*ۿ�
��;!����8����ݕ�!AE���|����'8�QJ(���)L �]�2ݞ~�Ç�L#t������׆s��z"[��/�b��q�u;�CQ0�$c�.�lc�JFTv�a{y�$k�G}�R���E�����B{�z����T)6K�5,J ��V��1?�`b(��~�RlS��s��m��T��+����;��o�ȑ��~���mo�ּ�nk�@}�4Yh��Cь� ��̋0,���#��n���H�A灇e\�2 );��Z��cR
���^/{���B��f�E�܅a�� .����$I�ƺ�6٭�S꯭�� K�%;�OӢ3�����c��f��M�;��
�%+�(���O{�ʲ�M Ec���􄏇
����:iĶ97u�<��G~�"C��ɋ���$x@5
dl��΁�Qd�C�;,��n-�|c���۫����2�:�K���B8�.�����9���	Q��^����@}׭uZk<����J3��]Y�/� 	�©2|�g�G�%�{�����﵎M��(��E���V���HH��CzT�+�9�a�������`1k�rF���Kq!WC<���m�2YE9=&BNs��f&�B�c��v0���4@(�����g||�B̔U;$�x��*Cܿ��_a�K��.��OY�#�D�v.����<�3[�%1e�ȅe�in���X�;$��f|�:dZ?]Z>ڼ�4�=�p�����?�qB�6O(���Z�-!�r�=O� �d[�V��[l���L]���oH�֛[F�;�i����}삯�7"�i��BY�,%��W��d�X'��brm�(���|�����+f��5Usj���m�yu�`�i���H��׾�cl� ������M�"v�i��L�^�Nc�%�u��ʡ�'9�F^����j�"��-x.:�2:{u�Y�8���y�/I��R,pkrE^!:[���^g]� �2��J��C7u��Yz���!�< w�j�߸˭1�n�j"D�M��|v.���ɲ�-6��h�:����O��	�v,����q�l�'�n��ٚ�+uAb@�@@�~�騮˂��r�\���,�R�Y�^�)�/��K�55.b�� ��+�	<���_�*W/7�*X�ez�\��1�@"��9�{ �v-ee;~�¤$��!���|sҙ&@���7R*E*�0�`	�ͅ�P�۫�2��;ma�+[G�k�p[��(�_bRYg�<��odCot�G��9��n���/;�|���i��ò�?����QT|�C���H��>�X�s+Vr��G�T�[+�3e'Sit�����"j�v�/���GA�kX��k��u
y�Y �t��������,�kV-���_��*̚�{��TAR��y��Q/�����7ۓ�s����*k���e��Q1k:tia[ݗ)��X�S��h>�n]�V��#\P޾�A�a8wܣ��[��#Lq;�I�UX�#o�e�n2���C��K��p�T�Z�[�L�!�)F�������g�}N�&*���w����t��"i����t!�z}#���ٍ��WO�*Q*O��=��s���˯k%T�ĳ�E��z�w�T�שͪ�N���4���7�i�<<�+�����-v2�Z�4�f �K ��7M�DN��<Ox0����І(ѱSi�xɤ�9,��iG����'hT� �N��K��a����	��幼�F���� %yV��h�P���y�zA��
�;i���rD�W�4l��Jk�e\�qϹ�p���z�&�IA]�RW�uA����g�A,�E��}n���S�'��=t���/gF�%�H�<��E��A��P���Yw0����spx\���h���M��Y�0ld1]2ѓ�]������~�⶛��G|�[�K"�����~��Թ�t��B�dD�cą�u�/sy��Dg��=nxL�c5G�7�ݕ�A5�yI��n��rF�	�ۓA�7��>|�����~�%����zI�8�߁Ow��کO'Ī� &���y�`�`j=�5���c�몮@evČ	�gY��v�a�{,S��I��g`N�bSa��?�ש�^g6DGȌN�{���Z7�"�.T��'���O�b_�i�1�����Dr��au�" ۰�@4���mZ(P�w�6���$��ݞ���zr��
�1�Nh���h�MF�bN]2���%���HqL�m���s�e'7�e�����#r܁�%�].�lx^��n���R��>t�4ox}��Vw��T����\�9�e_O�s"���]� )7��W�u����Pb�x�Q1���4�nTv׳^r#�.�lq�~x8)R|�����I3/Hq�Ͳ]E)�1�KXW5�@�-��j�ΨV^��^�܈��ݒ���ٲ<��HIou�L��O�@�Q�
Üq��^�4�\�;�yr+2�4���9s�0�����'| �@Q(�u$����Ըk	���M����`IgS��%��k�s�@\�q��Z/ݙ�1.�[?�6��T�DQ"2?�b�YHÕ�O�;��[o����&+K��0dFe��C~|~�� w��&H2�e��TÏ���t�/j!4���&�-@c"ej>������ƈ6�7�Սk��f���k�-���w!`O�?V��@~�R����E'��,�FFmu��8��1���@B�즁BıJ��e���z���nS�9O=����2�p��$�\�-�*V�4j�t��_ o��`��Z]���a�OZ�:�����b�������.	���Pz��	�Tv���z�������N���z�eu_� ȶ�'%�qJgV����t�\����U#�0����T���*����uA(	�W�I@�N���Q�D�n�>(���vK90�8��E�
 Q�S��!�|�!eՃ��8(lG�_���_d��{�����0�hnA`�_����"�m#���k'�Н:��م�Y�TE�]7�^'�;K17�'��PM��z���D@�j�e��n��ݑ����i���n"zp��Z���0�OFǻ�8-(�O׿r�B�V��U<��g?����J����֥9o��5H��ct$�y�����b�|ΑA���j��)���a��\
�ױ�y��Ɖ��u�h�X��j�`��&��
kmr��ſ�ˋڸ��X��ݣ�-�R�F��"��?W\A���5���;����Y�
�3U'"���*Y��!���X���m`��X[HhR���
�W6��-5�S����=�1�Hć�����ڸ��^�B�����ӂ=�ASVPI�Wz0C� ���1ӈVn�ai�۔�6���T?�������9��D�B@�������M���{G�Bx��
|hs�0�I��^�2�M��ZZ0G�R+~]�������6D���qY���⊛�E!�gP�9N�d֘4T�r���w��
�����B6� ?�U���V~=��tP�w�I�ng��F����D��5�P"i�QMΡ̪�G`�J�M=��1��?�������M��o)C3�����d�nb*
�y#��(iU����k���{`׬=�B����X�ě��L9�~p�����'c�(���]F�}f��S6R�" q���4ͺ�?��p*Z/o�E8�C�_�Q�*�Θ �̣D�E�#���4��̏�&�f�·T}Lr*���A�Ud��T�yUw-i�2�33��>)�M��`?��К��F_F¡8o7���ȵ-R�:�%���Z��5�t�S�p�>h��|,K�_T�J��Q��{�H�'���AH�at��r��;KjgE��g8��@۠������W1��b�Cd9�@/���A�)����$�:�L��)�Y�8�T�cs�lprR���D���y|����S��t�&h���F&�i���i��bv!�����F�r�y8�E#y�3�k^c0��\0�rU.Ƌ��-�F�3�}L�Bj�<(�ު7Gx8�'hi�fb( {� vg�{�C3��d^m�jw��G�u�A�Xw��~� ZlF���
6+f\�k���99TEƠ���!_�%`�
�y�����abI���6%�&�8�!.��4��Ep�=��8�wv�;D��ߒ�����Q5�_���(�Xç&�8
1����3��n���{��p�쏩g+����������N�v��yL���Z�7�F5iE<��)�+�PE�uk����� �����G��閲�N?_�}lCd��ۗ��2t�b�:\řj%2	;|[c��,��x%�5�A2i�=WvD1�K�C-� J�/G���K�v��Oy��D�2U0�\��T���:r7���F�L���Č7}��-0ZM���En��Eu�r���7K��*���KБm�څ�������,��3�Ÿ r�9x�����!�/%Y�#��u5��.��ff�O���Ya6�L�3-���~�(EX�B&i��9bۜ��G~��.ɑdI8�S�4�'H�q�\���K�h�`�\�0�HS} =�|����9ޱ����da(�Y��5hH}yn*��E3����0��q�g���l��;�_8&��X0[�ߴ@�6Nq�e�V���!rh����>85��]�S�c����ɼ��9��/<���&�G�޵��?�^r�edJ��kyf�Q�X�K���|Qb���C���I�~�Dq�8��n����ܟ��M��D]Jҍ6z�m�!�)T��H�8�w������8d^b;�}o+r�%;F��݆0��
C�T7]o����f-*#l��^{
B
�P��6�V|}r���j��T�P���k{my����n�9�9d�u@��Y�@X�(l�K���kz�#��u{�a���]E����_��J�+Ua���R�4�B�=�����\msPbq�W#XefAs^=��>K�Z78��Q�~�.N�X�Q��ǉxC����T�Y�K�K{f(��k��}\V?ΐ���&<t��9��F0�����PH�,w&P
?��Æ����υ#�B>�#�e6է�:Em���Rƣ�;��i��{�~�������M�2<s2�����K�C�������Ƅ.�l����b�t㮁������,j�t�
H	�'�h<�:���qA̛�'�z�?@�`@���@����T��4���|�@�b�����)���y�`4X�aS���$��5ʁ�'�'ٗ&����n��΃�>�f�Sx�;�J1�+ӏl�5  �fTOn#:٪Q{ܲl�	Տ]�F�}G�{�_�N�%#���a?�%�G���Lɡs�3�(&?�l����W�z'�^���0�
vj6Z�)��yXk;auC����vBmƍ�1x	�xhVv�c;���p��A	�5`�y�N��ӮZy^=�xT�N4�PQ�Ѩc�@���U��n�۱\�Tk�t�����e��ď��i�,/X��+]g+�㹆����J�R�R�7�dW}�ڵ8R�N*��$�es�q �=��2��w����̏bd�#�|�DO	+�tC�Y@�`���T@�P,8�6~��?�)4 _��	0���裷j���=�Q�aO�O_g�yǏn�C�~Gi�`���1�C��
�9~Wd��\��v!���P��`'��}�c���aT�	�t��G�,2�"YLZ���{G���ڿ���/;1^/�0����Z��=��v�p����r��4��(kn�{�9�����X�h>�,� Ȑ4�O���s��D�����m��j���
Ԓ�DSW������5ȼ-�|�H5B��T�Z6C#:<5V׏�I���\q�!r��`UO�C� E��NB3TK2u�NЬ���9'G����c/�1@�K��W;�ƻ�qcd��#�?u2;^�i��*ә �<{��㮌
.͍���TQҊ"�`���Z�+?&��류�9~S��H��|�>oR�:(�� o5���8�C�n�^�~��C\��{D��lxW/�Ƶ��	x�/$�1�Y�@�vk��R����U}������I����]14t���&�&r�VA4�D���m硚� Ҭ���2�	�I����8ڦ�bl�����ε�g�P/e}�b��!��s���c�J��a<��e�+�:��f�]���JNp��m#��m�W@�"ĤZ���Xɫ,��.��W�G�~Db��K;7���nK.�nS0���n�r��J˽D���T�������9g����i��TM�mYN��IJ��h�x8�����\�	�� �m�5�������Q��4��@�t|�d���q�@�
�J��-�s������Ӟs�!k�+�T)�!�!�D+���Q- ��yr<iv(��|"��&Y����qƜ%��5��K�H�uȢ0�T��b�#}�M���[�Cm�tO ��;���3��A���-��B�E��]:�lH
l:�'��@�@59��'�z���/m:�x�K�+w�8�\чymd��%RXyD��$��s
,"�v����5�rܑ-!38d�1�~s��m���,ˡ���3Vk�6�/5�;U����$�>����O*~�Fݳ%���:S1J#^fSh�L׎���g����p�N��WU�2/7w؊�lU�b������5ZW�{�+����d���pEfny�Gݐ��d���ya%�7ϑFf
(�u�l�s�9$�L�{���i�va�� q�=�_H�C��x)l=G,���-++��?;�)�r6n�14��(����̐���=�vi���CAP`�~ލ��y��罍��q��{�o��D�!�k�tl�eC�D�i�p��n�q筲I�l�[ʱ1�>?t��pX�8�*�`�9���m�"���9J��32����y�ш-�Ӗ˙����jU�e���E0�i40�vu*hY�LL��.�\/�s*6��!����L�V ��-v	�ҁb�{�N�̚s��m>�kt�խ��ɘT��}��[鼠ݚM��.��w�<��ԫ�S�5:>PwO��uٖH�y��| ui|�ş(�4v�0�+ ��E �p���Y���~�b�w��|���B���Ԡ��zte�B�6�kw-.i�wYM���9Qh ٫s��S�:�a�'��@�E۬?�G�7i��G�q£�&��4a��q_�CF����&w hc{�������$�o]el���[LK�`z	&�/<�.�}r����- d�ׯ4]��Lb�0JR�}ޙ�>��i^�Վb|�����3�� �>��W�}k|���.G�2]�$�4v�qXI��s���GE��AI��O��0�߇[/��*��G��!D��V�W�·;��~Z��	g� ��gՊe/EM�ٲ>��Oh�H�����n�b��Y���V(*��?4�f�s��^y�6��0���>�����ĩ�V��_;n�<�S����ĽRt5+el2鯭 �"����aI�4wq>"�b7��F�������(�����R�S9�ʚ�oY\iA@�o���1l��W��'���Q�8��9!��B*{8u��MltO'�|���.E�IT
hR\}�nw�D�_3��)H,6�'���vB,�Ff�f��DB��\�L�z���s��1&������&#["-��k�lN&�0�J^9�غ��[����871�:�G������)�D���Y0���<�h�ݤ�FS��ᔑn�B/C��{ǃ-z9�����u���������<D�z�K؝-y�i�ryC����������s#���/n�u����鍏^y�DSE�����Z��f���!�,x�L!ƛ�7*Y�E�:�������`2���(�7`(��l�gk����^�a�B������ҘC0^5I�x:�s��ΰ���	�j�K�_�f�������G��[gs"p�CWn"�ש��e�~Y��(�
R>�X�jșL&eD]���Ked������c���GC�o�$�����"�ྮ@��ؠv{yTB?�5/���p܆��ʋ܈F//�ܖ$�\3���Ƭ�Nxl�!�Q\������ab��u�r��:�!^�N\���_;���G�p��=k쎝K=�>GqQ�(X��
$� �B��I�dC���4�ɣ��DJ������2\�0� iN�z]C�O�/hV`�,��_Zi����X�h�Y��~�8��6)E.�l������zJ͒�ƴ+f�4̗����q.BI\�*���UxN)��a�&�<+���z��t��K8���h_��W�PR�ǝ�վ$�`�]�0B�����σ۳�������Ph�&٥o���P�s��ʳ��V\L�LA$�a$���p�1č?���Hn��'���ڬ�T�ӗf,��oEyM�C��='�vl��_�۰���o( �\#ф���[�NW�J�{����i��%���lX=�;H4�ږ*I<�	kC�3L�,�x\�A8�6�0�!���G����TM�������aX�6��L郯TYr&�'�|#]r*����l�y�4��K�ӱ�2/U������@>6#x%�[�ܲ�Z�ov[��p�:�̭�M�8�G�:��i�{��|q�܎K~�x�@� {�����ߐ�\Y:�{�`#8̾|>%���H� ����m�w�m���k-���{{h���}�Y�J�̧㫁��� ��Y�N�+��T��)��q~3Y�Ĭk�*�	�܊���6U)�mO�ɣ�H���Va�0&3KR�J���"/[ҋ�7�l�	�?ĥy?3J���F2��"]8dvo��h�X��4�
��_.�����=����,x_r�Qs��S��\I2̻"y+�n���)�����̡_��u����>KT_�wgK��X32�l�yv����a<�;I�i���֎43��L:��i��4��ژ�v.���B�Ն[	d�J(�����ԣ~�+*����&�T����T����[�(_-@�9�qX�iX�ܞ��Ym;��M��A�Ƥ��O,���$?��y��4`	~2J�u��X���y]{�s�HlҴPߑc	��]E9E����u�����UQۘN\7�z��v�вJ\��	4lc��-��m�c%��JP�dC��
+A�[��(�����y��n ,�ʼ���Z�F�P�M����L��T���d�5��׍���K��xV�K1 r��00�!��0�"=���:_�T���.�N��@Qok9pk��
[0'�PFLcW�sj�S;e*f��2;�#;� ���ZzPxۦ�s����:��#<��+m:ܭZ�ສ|��d����gp%�3���|�ⷄ��!q��8]�}s߽�2Wj**<4�dC8���O��%B���f
��ͯ�r �'��?L	�=���
��PsN�H^�}q)	���q+��e�m�䰞��C�+m���/�(��|�Jfo���B��a��/P=�~�t(������|�ņ<�Z�^g�b[��I�oԫs#p��+ȭ�[尥qra�;c��K�WiF0�P��~���&=!��<Β�/�[/O�~��F	<���g�ĩs(��*b�4��O����L�����^B(w�b�N��q�
Ł�L^HEE�ʼ�D�3Vx�d�m�Yk�C8�|�+�5���9��������{AVGK�s��}`�R�C"�#�a��>�!?|mC-W����:��1Cu�'~�ԙBq��N���1,Þ-��@ʞ3�mrA��S��ɀw
7G`n�ɇa�ml�jK��*R���e�˦?�i��Ĵ�q���_YUub�o0�^ڽQj)��WC{��K��p�_Æ�S����\�rh�uX@O��Z��_0����	&0�����l��@����DsJ|�K����(ߢ	3i�����̷�3g�c�x�n�(�ImI��I��/4���3��ƹ���{�8��	�Hy���L�EA�as�}S�W�
gw�U�1+�j�����Q�L�*uB2͞�X3����(�!J�S�f���w j��P'�A �e�J�FC�ȹ�����Egn;D���<k���I��Eg!~�Y�ި DS��8����W�-nԱ70��g��H���$���)�(7�r���^�#�.�$4��yx5�(Jz��a�c�Ghե^6�=@Y���=�nǬ�Ʉ��੦�knC'y��Xh���:�~�OH�t�]?�E�H�|W�-�~�f�Z�͞��*x�T�dj�_�1ߏ5STI�M�� ���*��o�ü_��h?1��#5}�d<�ۜX=�oV8��h���Q`p��I��F	t8gZ�n.��/$|��Ǝ�^����O�L��+"S_G:�0�3&c��c�f�EP�ۏ�Z�iD��c'��M}�3{H��G�I�Ϟ�������$�$�5-+a�ǃ���_��A�Z�%��G&��ǌ�z>�p޹3E񦻌�K���2��i���8�5�)ĎZTm��M��I��o=1���e����2���:B����WkR��9���諐���d���� �"�*�V��D��I����W/[]��J����Ϥ�o!\������\������K�[��-�	}7Lƅ{[0Fe͉w-[���4��a�Zg�3Z���z���y6������Ē��P��̛��h���&�W¾�l�iqd���͍Ȉ��_�yt1�氼|f�vj{�6_�y���)�Nm�J|�.�z�	��Uх��T/n�n�%$���	Oz����k!�ϻh��jL�=0'�����)��z��:%�0��?�)HZ5@�7�p�bp�X;�[k�z��d�^^c�f�e)4#��~G�a,�#G��$�%�S���|���0��P�X��)��R��2��%�q:� �4��15h4��.:Nυ�>���yϭ2�x~�~I�XK�Y�=�
n�	���02����*g�������vN�itm��.� �<5EiNes����`zE.�7�N3�����c��~��-����˹^���9�jD&�#��	?�W��;k,O�Pqی�Ya1�J�g�u(!��s:CZTܺ�=Bx���Rc2y�j���.�� i4Ѯ�����h+s�Q�|17�YgR�ao�)�\����M&����#𝾣ϗ�wd:�5��潯g�;)�:���<Бa������ę��:<���%+��b�/T�.�Y����՜�e�����9@�*����uc���ra�ۺs���ޯ�;}���@
0�� �C0��F�Ț!��I�}�s�A��m��@��w���&���Q2�⦁��_��F�d��|E?��?�S�,7p4�b��RX�J*52���WD�Pr1:�Q�c~��n�{~�9�۴�&���1�j��$�q�yx	<�)l;zc�${�)R�k˩Z�M���y\EM�A�<WX W����O�v:Ƃ��(�-|���_�U6�շB��sC�N�6�@8+���/��9§�1!:��`�V�f����}�d+ʉ��a�&�v;��ϻv���K�'��υ��U�6���̧��^�aa֯zB�Z�����7�����a~7PnI������\-�{��y���R����){�	_t�M�d��>�~dS�ǧY6�p��P���4g���L�� �R�P�6�{�n� �4
~cޝ�Rb1!.�gv�{�`bh�!�l�Oe7�I2+6p�t��1�t�����66 �8��3�X��vo�S�ې �KMh�SYaI���&&�peģjY]�>�~pv��RaIG���6[�{��W�0��5ٕ���5�\�w;o��ׁ`-���@~[�&Q��b�cV#�{�#.&8�a����T~��3�BI��'arVy�턬��ěm:�#���h&���|����G�0��B gČ�>�6�kAhW6y7��ˎJqU�ы±�b\y&��\(�O!� B��Jz���sҎ�r���Xy
g��o}R���]��o���s/�
�Iq�$>�cԮV]��>Y{�Ȫb���r��Lu����YF�Ry(x��\��2�<(�����2�.���u�WEm������g�!������j���I�`Eט��:��	���i�~�WR��~SJɮ���	/�s����A�{��L� ��լ��rm��r1���8�epyi|o�Zz�8c�(����Ck�[z �@.�=�Z��}z����n�g�A�r!��'t�l>�:[G�%Y'a߽������H��,e���V�I�`�a� 
G��9nErGxO��D���"�5���MFF�<i.��!ZQ�}~F�x���S�&9�-YUd����e�`mi���~(�������˱�,L?�a�{�$u�Afl�,΀f�H��K���?7������֊��(��<��(4?gT3l�d��1��@��J��љ��#�SP�	�$�Z����E��/F���%^�3�7�hZ������A&��Mr��w�:�M���������у����[@�C��$pvM�ID 8��ɠ�f���+�y�i�ۿy���hG>�S�33VYi�����1�P  5cҊ$V��>3��ɏn�F6�VO*��F!�j= ���I��.v8�(�	�BAc�+��DV�!.O�m��ۓYoh�ϛF�Bd���A�HX�m&�\oQ9�zr�M4���d�������Ux5bC�Ω�Gy'���Ia�b8��!JtVB,0@G@�5Zz5���BݧҚ�Y�i��b֍n�F��Ж�%���ݽ�4w�����ԣ�Ϳ�1e�`W���%2��Ӣ�x-�Q,���|�t�G��5y%��|Y��G�r���s�ܮ��@E�V���V!�cp-���da��T<�/�R�3}i�ȸ�d9���L5%�0ϱI�����"�)���r��	NV�Fs-u:��K��|Y��������&V����9�@~�jA��|)$��;W�������~!��K��)�'6�9l#%�'�#I���B>C�ug���g���6�{�����f�d�`#k��6�1a�Qg*[cԘ8ьe�@h=[c�'�FiB�!����4:������E�h��#dF!Ǩ�
e^�:D�8kT/8X�]����y��x�s�3,膯���y�< �|?�D{u\�'Y8ID�<��ݧMv צ�g�Oޒ��EPCs+��D~��e>��o�(��ႉLȠ�{��)������[�i3�B�lN�Q3/����IqP!���y��a�3��Ú3��khk2�V�S��O,3�b�4������h]bǍ��ؒ XI�
�X�I�t����������7����R�;[!��'f���?A��s��GO4�H��"O � L��̠ "����m�ً$Ū�A@rڗ��=�?N_�ro�?���\G���Y:$[9�j0;����t���54�P}�q������:ǿ�GX�VN�kG��>?�)��E�D�p��X�q���:���O�O����T�wW`���!q�����4yB�D�ҳu�w����Y=t7��i��~�'��fs�����x]���.PS���3m�gDf�ݛ9�w�i���"M�Q��1BDE��t"W �E�d��_��ڎ(j�{N��Y�ֵ��K���)����[;f�M?	N2Xg����r���bq�T�I����b;d��=�8p�Ϝs��4Y�tF����6���a�-�]p�MD[��߅l[��X�zX�pؽ�lb�UX��H��7 ��}�E���9����$8�$�
1Α������w��3�O� &��#҄��X�^��6��F�%�-ʔ���c�T���R�ad�i!��x�K��C�7�	�0�����՟���{�O &��)��>IL�h2-.�I���!��E�wSN;��f�
<qe���xK'�x��2b�Y I�N�MM��}��y�����;����r�9��>Y�v6�a��/.K���j�_3붣�靁�t�W��nH�z��fqy��%M��Ӊ域6�v³E|*Hm]�\�22�fG�f�X+�o�z���&b�Fً	E�ʨ���4��{�=W�2V��\XelQ�aM-?9��J]P�@��T�}�����a�,���m��D�T��Q~t6�wr�b<����r�J8T�N~`�>�v��;��Wt��m�J�9�Z�-�7�
�8�(f�R��e9�h]:O�Wt��7)�����ܠ�D�������42ySbP� �|��@�6x/�8w�l_���gM�-#0��P0�x��罥ܾ=M�3=��#E�����Ń�mf�[3�u���qeK��S�h�p���^V-����\R�[K5偞#��{����뙓���$�P,W�e�މ�5��E��T�W�O�8���dp��YQ=��r�ai*w_�_��U�'ժ�9�~;b���I����B���>�L쁋��Sj�������WJ�kJB�� ���4�3RT��;Y��i�P�u�g��z؋[�����8���USψG%:V^�M��v�2��#�R+x��l&�==���v��!e^���qo�Ng8��n��1�͓��=hM��Ǜ��vw·b�w��|�b�\uT�u�d�i�b
��Z���J�BJ:Mt�~	PI)���k!U�ӡg՞��
9�~�XՆ��s��*�'��&�_�`�%��R�(�,��M�^��B�*����������h'��u?5	�%lb��%	�,��Bk�M��.�������|�Ó-x	\6	�O#����X�+Q��~4o����	�`㩞ă�LG�=�˸��7�E����[$�F_����/wvg�~9�e��b<�۸������pa����8&{���NIa^C�����K*��%Jrt�,`o _|���B�x��./�,�E�X *쵫�N���e,3�QC�A�`�WU�8R�#�R#��ܐCܔO"D�򣌟6�U�&l�!_,A!��<AJFAn��推m;���L�1��l���E}��\��+�w�qs���I��d��ǥēm�h	�&��-��{|�f*���/e��e\��4���+���5�A0C�_�䣐���F7o7��+��ǩ�߭���G047��I�»5%�D�����oE���gTW��=�����0��F�	����S��'�j��*�n�v���W+?�F"�H��y�Z ���׊���3Q��e/���-��OX$�**�6�ϥ��v�uC��c�UAJ�a�t��&hk��5��, E����cXo!�C�p�A6g�Pɔ�k����ő
f�<(��B�3AT�S'Q�=��<9h2A���>���;�X�Bo�����m�V�IZ�s}eb�n[iz
ʟ">Px���#��85r��#��PT�Exq��4�g�=گ�i�m+נN��#��=�8��-^�,����Ԥ�@}�#�R�L��t���/7���16su�L����J.��6/�}j��V����\��l��W��7U(|���"��T=x��<�*2����xv��V��H��K5�uք�����L�d��v��Y�5WɦK����N�:�6����l��ظ7xO�в�<�<<!'?o�
F5��l���>ј���a�l�v�vX��HbՄ��aF!�F�_V��^�n�dS/YIH*9�Q3!mb^��@hP�4ڄ`�'�BO�?��HbQ�5Ү�R�k�l�;���c�YV��rvc��+��q덨�ʕ��ŢS�d�p��O�)�]���u*ѵ�}l��W}�6L�rq�˸�\��/ �$)�H�6w���τD^�S?�]���3�
���*z_~�U�o���L���4�e{r����]�G���~������x�$���Wk����(���V���T��9iG��=�wG��C��U��1��Љ�2/N�L�]�'���IZ��)ʭC�0�n�?�;k,���:�×��G�y�dN��M*V�:ӗ��1��-d���L�7"���z��W	�+�H|��8�]��9��߯/��G�4��)��$'H�NHq��oP�E����\|�0��$��D�WT}ԑ�W���ef�i.Ln=
����3K�JV6�]%�B�=s���y���o)R��Ǿ��X�n�Xr{�8��BSc�Q0����3�`�Ngj�7ŝ^tA��n)�
��3�Z�z�e���Y�r��&�)~�fƮ�Nt���i��s��o�.8ȄMSU1%��.�����b.OL=�Md��uY�ݛ`�z�D�q��ap�+0O��m�_?���"(A�@OS�ƴ[��x���>���a�/��	�p���[�^�yd�����n�_iܐ��3<�=BDwgT���b+1>�f.��o�0���hh���$��DB���l4רW�V��	����/SW�ʛ��$�/9��Q&�MMvF>y�)�,ֹ����OEp��N�.р,��
�vq˴��>7�z�܂�J�͓�|]�K���@����:_<�n�]���6�@b�}�N��eT�K�`q�w׵	؄lˑ���ic���Iy�:�p�?�W+�T)j�@����;�(n�b�:��
��pʒZW���/1��ВL��:a��.���f�Β��Ɠ�A7D���Z�Y~�ㄪǕ�PT���	AO�c���qE�n(��+��9(u,`dTG�{�6 `F/�+�+���^�_AP�v|�xA��#?��}�Rػp#.ۑ]	�
N��3G?�L���K�Ƥ�^�����>{�����9��Au%�µy���IW�)����V�C�yhd�w�P���F���W�tu�(*���#B���EN�bِ��:���zmTrΣ��Ab�i�U-DC�ג)��b�a�p�;��>&�e`J_�����0ȉ�Ic�#e
'h�?/��
m%	7��Y��x;��<A��V[��p�����]T�2���"i�d��� ia(�n��\l���s*8��^�L*��%D�X��e���aF����ʉ�y+��aH��܆"�L׻�s���l�'�h�?��I�F?��5�`6~c�^YE#���r��xHТ����i��T����1K���eg�C(�k��$j� &	���Z�Ny��J*���2�/v���Vs�6���o�٭����E�t�n�_��L$]�����l�������v���D$�u��W��9�[���s�C6�a����<c��C*h8��?�9��Z׸��U�u��8�}//��݋�`x�a��|#G�|X(�~�@���<��H�픹|��)y~C0)�M�C�~��<���D�V��6���C*��A�$O[ǎ�2n��L��>��S�S�i�	��N�N��A�c���M�͗u�m-��5^kdۼ�E�S�MU~<5�t�<g0�K�LAo�D�*�7Z�_�� �".s{Q6��Z�^��,d.�s�\x���=I���9	��/ѕA�h=X����f�p�ukK8}�Ծ��t�����@ۋ������cl-YU#G��d�$v�Ӌ�ȕV�*�:^F�0y'��)e���_ ��*�?�و�H�@b98*����A�w@k�n�c��(dG�D����f�]	yfKn���H^��o�us�ֈ�+$:U�����i�W��Gл�X�ٱ"��l����d���x�U�֝�݃��Ȟ6v!��ES�U�WC֖p�v�ԟ�%�ہ�	@k���$�j@QJ2F�GSu�Oj�kK�;}�ֶѽ�}�yzK��`c�~Ĕ_�5�dnRc���j3`aQ�_;�jNP-�+���� 셁H`��x�	`9k������ᓃh�����?٠QX��X�R�W�H���@O�R�*Ϝ����8o�HZ�s���V �U3�O�(�lUI�!mх�F&6T`��*)�У��퐭�h��ϛHt�)C)2�b îV��
gW� ՛�1�ٛ���R/+�'zf@���`�{�y�	�^�����MO���#w������v�1���Tvb��ۜK��p�~3I�����n��/Ѻ�T�B�w#q�%�`%k+���	Aj"�&�1�K�Q>�$&�Ż�|+B���.XϗT�>�D��nt�ۼG��G��l��1�;_��_}:΢7�����|P`�>$�E ��� ��� �Rޣ�+"1�X,���� Dm:�o%u�2�V�X��Lb��禍�0��s�q�^�Ι]�4�	z��qX'<\�xU�0��_�vnS`�˞�R�@��Y�F�����$T|5�\&P�h� ��P���|��q�;�X!]����<T[��z�g5���a�SA���n,������+ܾ�mts�,H4Ufҥ�
��H�KP�u��j�ZER��DKu(5@��hQ��L��i`d%��`{��c�%��ü��?��ӽ��,7��ww�w�4n��@~dGJegb�����#@�?�D���d�v�S��OJY�an4H��_�����ѕ���c���z�����=5V�KIlvli\�.E3V�dxd/�uN	f����� ]�X.4���V�cX�\с�K�ն6�l=�bi�/�(�{�U�ܙ �r�4��:B4-��x2�B�
j�ރ��(�ǯ�9s���L _�`i�����M���y�%w�nrT�I��'8G��ؘ�:l�F�.?�,U�߆'���݇�s�U����Ž��P]%�Jw�M}5d�<*�����E�w��eC8ͻr�*`�����1w�O�A�iX��Iv�qae\l�V�v�wf�e!���$H� �wJ։��v�(vX�V������d�f຿�9b�0)µ$������	���j��ƙ-Fp\�!����Uy�g�QvPJ���ͫN5g�wVr�dKb�\�\^%�GXޑ�#�İ&\E���,�!go�
��LO����b].�j�h����K�0{>P�E�^�]�0O�PjS� ��F��I%��_�� �콬vZ��<DZ�J/����Oi2��*�[��(��ٱ�}���Ȭw_F]h��RCZH�
}�{�����vn�2���hJyx��������u��]3w�1�AT��s����'�:���I�첉��[�D��[|o
�w��ՁW����ȇä{�Ў�ES7�^m
k? �ֲ�g�'�;EN����-��w4ɮ�k"f�L�7��̐Y�?�,$1�����R&L���C�D���9��"L9�z���yG�B�4>a�Ws�*,���NLp��ZĽL9���ܞ;xS�b��8�SǪmN@��ˎX�4~�e�
����!@�#i9������
����02x��M^�����C&�H�Gc�Zi�Q���W�h�C��cV?�������E��к��#�x�9}jd�ُP�o�q�%�U�\BD �*�;��c�=�6R"�6�OR�Ȧ��n�ϑ~a��_�(�*�ʤ?ߏ�K��q�Ș�*e�`��\Y�#)VYVa�f�;����J,��dc���J
����*�01��t�7n���-��r�������x���HL�n�&��7�Vֿ���n��;د���2ҙ�7�L�-��X�i�0�߶f R�@ư�ˏ��)�2��$��Mp:~m��X�]o��q��}�@�S��}h��4�#�9�`��8$��O�g�xkhl����^���n,��7K�$����?,��(
b_�M�d�ʋ�؍yJ�8q݀\�^�nN����C�%�V�����$E�zv��N�=�xڟ���wm�Jo����b�;hlCY�,F��j5 �~�=�n&f\R<�+�_��?��?G^O��� 	��OP{���˭)����yQ��&x�]w�[�?$�{���svN�rx AIIk4����h�-�T�-�LRqK�V�-�n���^�����'p����KzP�2�n���n�5�}�H�o�.�s	Gi�eX7��]$[|a���Zܰ�
�,r7Q���H�~��T�*O�U0]���=�Q�,��M,>��as��7�L��2^������ڧ}~ƸӸ����6�b�i�Yiٓ�+�:l���T�;$��*ci���� ������-����4Np��>l�D����/��m��͗kB��O�9���^�X��>�2��8i��6>���iʹBR��!�E��������Y�d�.s#���Xî����E����z��Q��;���+���������׵���a[>�������8ZDy���r����4�,��M�e�/�=6��q�TNT��7�Y���/=�e���K��tߖ�:��p;5s6雂�����2��7¸�z�=�W�ˤ�b�%�!���<US�͉����,0�e?ĬP��ۑc�z4sͮvy�JHY�/x��Yܽ&�g����cH*����.�V���oW/����3�U�U��C�dj�A��)�tL��m���l��������Sٗ�h@����=�D���k;��k��Q4�=��YL/�)7DZ�i\��DLN�G�],���N���딘��1� E��%1m��^���3F�ܳf%G��$��K|e��?�E�&:g�䙪�"��'�Em3����s�z��6�K/Ls��񄥍C����Yw�?��L1�/���^���z�Z�!%dX}��2��q[���Þ_����;Z��A�q���^�Q����4����S\����!i�<���<]&��e*��F��e�@aHk�S��]	�c�������Pv�!��8�|"'�r����vH@� �x��!z3������&l7%S�̣�,H���@�-ښ�Q&�)s�z��DJ���8�YAH�u�?H�w��i�Ͻ���y�9\o����bk��u1D�2`������BQ��R�)vώ�E�I���(
�|V���v'(BYu��q����'o︠؇N��{����*���
M��H<��o�t�܎d:�ҼNQ2`�x���[Z����пc0U�QdE��n��F_�0��*Xpv�H��0!�Mg׹�at�[�$��{s���<��N+0m��h�N�xZ$FYϓH�ѣ|Sm������Of)۬<)��0�E�(����Ή�䟘�	W���R��Ly-穓ݗ-�fUJ�.�4��0����; j:�ã@D��!�����L���bP�I������LD#��ES�Gd�u {��2�g���x�)���Y�ݜ15ҿ�]:I��V�"%�س-���1��-���Q�E��Ik��4�5�JA/��lcWWIдi��fr��~u���#5C]+6DI�����祖����Ȧm��@7a�j#�������A�Up���&-XֵZ��	����2;�H���@����cw=�}�&#I�c7¿��5
 �vUpa$�5��sv\�7M�m�����2��@��;L���H�Pj����U�w}eS9<Ng�c-MC^�U][�7�1�,��n���+�!-�x~�_���h�7�*��~���tK=���U��l�_��w��9��P�����> \���&s��-�Ho�=�ժe�O=���;�²a]�n���Y!IC�����#��L��/�w|�F�UoX��zZ���D���3?�Dt�(����('>��gL}bm�Nz�^�:��`��׵Ś��>�B�(�+��{��0��	��`h'BHu�J%p��q�1����8ܧ��6�1ڴWi�CҦ�ɎȀ�?�A�3_4�c��q����H���[��1��!:C���#XV���3����- o;<-�*�������l��� x-'n�i(ڵ3���o]�~x��t[�oe�+6�{>�.�&D�[*oh���t�z��ȵ��)��ւ!Y��o���KM0�pS��mͧhg����.�
�C9�e(#����r��x���[g�* c�|)�H��>{l$����<�z}c'D��b:w�)����#r7�|���R^����V;}<�wq�v�6��ٮ���!@j�*F�0��g���1Ǣ��o����
��B
�C���ʆo�����[�[:�6��L��U��2�kQ9	?٭T��v4cŉ����?���[�����i�xSF)�xy<v�6�ed
'���\p��*��W�J���KwW�#�%i=,�I�uRT�;(� -]w��V��H�,�:a�_��.�懧.:pO1����7���h�VG�
&e�1�FLe����:g�D94���|��-�������T/��n!}�� DX����j���o�H����_�A@�h��(rlH��!e�r��]Y���^��H�����O��]$�6(��@�n�t���?�u�Υ�^1�ʀ�}>��	Bh��H�?LmY�����f+�=Q5V�ίٮ�)���rR{��=�Z����R�LUWh�k������)��e%��ʠ^ן�n1����������]��x`��%GBD0���EB�}���g�Q����=��IY\��HIQ�4��hr�L��ϳ���S���:Y@�=�nM�
	 ^EkB~��=��p��<Yy����}�xd�}pE㣱Ր#R@�h��R��iӹ2-[��~�0���b����\�F���AҘk5H�]�k�ʆ��5pW�@���E��I�w�}��,j� �z�W���T��={��0~R��ܛ���8��6�˩� aH?��;�\��,&Z.``87���q|�(."!��j�&u�0i�xA1}+�]�+ׁ+Vg�P��!3K1!�ȹ�8��굴��M~�f�t�+��~�q�!ڬ�پ8���Q�[�(�%U�,���4������Uqv����5���4� eF^��8鵱� ڿ��#��c�@�d*.ЊܲȺc�Sd�P�.��������ծ8���`{~�+����Ѥx(�E'Z�E��Uߝ�w�E����q%c�{������Z���]���"���"'��!|�3�� eV!A6�g����g��o��2�ȵY�vz7�䣟�����Q��Ty袃�JvQ�&^��xdro�٦}��$�W0GV�U$䣛[���F�i^�������6k�ޭ�\W��I��6��U�꨼�{̖U^c2z1�#v�2o��;Y���qHS�������������^��^{J�(��/�խf��7�3R����ry]��F�@�6��Q��_���&k���ogH Ƚ1�p����%8��X�?�]�t��R�h��V���~�=��G-�J�����"I���s�(d,6D]&�2C��GI��џZ�+�$M
����s�1��yR�(6B/c�9��7�������t��[����w�ލ�
^��S���@G�c�R���{ه�n��)C]_C,6�|m����EU �h%0�����;�(��כl�&�R��*�H�ܢ��6�LՆ�r���c�1�;�q���W�C�f"���O�l�T4�j��j"M�q���V�Q�U�Cӻ�k���9;c�07֜%�/d�ˑK�Q�n��_̽(v��[?)���7{��Jð���q�|��;����L��pZؠ-�����������]�f8�w��;��$��"�^�<�������dƂ���8c�%f�ĆM�Y~�EFм,�vg�qɥ��T|��8� u�>7�q���U��Bd�F���-�Z�QSC�ھ�$�PjhFT7@�]�"���76�(M�0�w��b�d�g����u�D΁�.���X+����7�c+�F?�R���˵Epe��p<�U��^�KuE�z�k��s�G�P�~�.{��Ze���������a[L��ѷ�ٽj�Aֽ��<{y+a�\
9 �d�''\0�YE$(/�G���*v�h��6|Awx��_�r�佚���U<<k/��
�/!��jE,�G�͟�u�߇���
A������?٘�� E�	���R_�|����aB���Y��sv����.��c���#)�Z��ŶӉ�4 p�i%��~��<o
q8�r��<��X&����뺇Ϊ]}��eW��r��Mg��4)�rz]���+j��v酖��.�(�s�������In�b�����@*�Svu�A+�̱���_��P��|3\z\Hm�.CEw�ac���{3�M��v�>M�>����E�A�W"H�"�ER}B�T��`�4�֊s!��W<Jl���?��� �L����A�Sd׆�].�t��� ���I��, �\t#j�[�F�hs#�=mI�PI{��L_�4gK���a���S��6��@���G�4����~`Ĵ�� ��\��x�;V$8�j-���*��&��wjyn�L%��^�Fu���܎Nɭ�}"u��kД���2��.�����)���㥑R�^���drF^o$xY��\�~����\�cԄ�e��F�h<+֘O �a����5����D�=�C`ɔ�����w.n��[�^"�*$��NY�9orA>h�+�����_ ('Nc�e��R�����J4��a�!��!3L�snbF�g�br m��C�WEhȸ*Af�܃]WZ��6�Y�]Vd(g�v�:_\�+N
��l]�������cH=#�K��7��pT���������Tf�=�m���6�
�7����Wv}N�w�H|���0	��+H��AJ�X�����Uu�~���/O���EiQ�J��R`�G'W;�}3,��vg=��Y����o�;GٺogN]X%�br�����q�Kj�dS��[�(�?5�����C��#�/��.�:F�b¢�>@BK���ga�&��3	�u�	~��n��[Z��mR����R"!%�R�.��+ȭj�H��L4����s����������e������l��_*�`.*�A'dM�2	�]�`z<"�H�3sG�%� \hS��a�-нo"��T��:��5$�6�9Yʽ�D��^0��Yv_�42mS ��d�0���Aҝ����D�� �'�s0_�=D�̅���5-������P��:�IU��Y�a��d}	�Sz��Tqt8�e���$��_8C�������G{��0�2�׺z���X�r�GIiW���G�Nh{~���]#-�`n�~*���<`"-�3��H]5��֔���D(�z-.E1�v��������1ul䷎6w�����sY��	q{�C�E<�(����Ϟ�ַI���#ܮ�g��0�~|ɕ�ϥڝ�+���+��/���|~Κ�P�E��f>�" !�ek��M��Z��g�� =�Ja���F�;6 ����|�ܔ��<����'˜7;pVt���?jȽ+�!��Ư�^7(��F�8a�ź��:��jdؕ��s���qm��S�X��N�2��� ��C�#)<�@(A7�=h}v�.��+����y �'����huL�@�=|�m����!a]z�sx�?[�
;�"��ɮ�v�A���@�m���'gS5ʘ�N�Rn�v����н���L��Tόa�r۔Y�V��z Z������*�Lqz���|Pa�<�$g�t@[�����>4��̕��'��pK�j2$R��Fç�ͽS��}L�|�ם˺-O��I�\	�4#;��u_G�V>[��>�7J��3\���@��S��O*�+��N��� �M����f���~L��1"sm(�#涧�ӿX^%�*%+��K
Y��h^���}���,��T����H#���XSx�BX��+����a4 Y���3�J.DuG������hw�a��P�dhX;�����#��N���d"�4���!AK���0�ua(�/7���H7��/1�6��	�J���5�0b �a-��y��2u�]<��M����v�@B�,�)�9�R�p��'�(��X�H "n�WaZ�J0������&Ķ՘'�1f����g5�.�c1L#�ѻ�.�e����a��E.�w�!��H����|X,����Ĵѐ����C̃ �����*�Q	inzr�Ӊ�
^.����?�<��5�.���UH6���/��u�	�>;jF�_�R�a�$�r�o��r�d�`�z]}:��o�]%�g�9@ɴ5
d�i��p�B��eE/��v��ߢ�9|F�?��>�� �U����̌&s~[�I>����%�q "���ĿjM�6�r��(�H-O����b"w{�x��ۦ�M�\7������(���=���2�t����#��N�1��/�7$�-N(>��y� ���]���ML �$KAf��gYq��Rm��\
��*�U� ?�Ŭ�AU�P�L�`b����> �#�t�4�t����0���3+��
�<������Y�#4�M�	�,n ��V}��<�"�������0�m���\1.ipT	�6���T��o�#s�No�L�Auy�5�������S���M��R ��e���R�z
fy��%7�+����#��g:t���Z~�K0��Č�~��5�����㶪�(Z�Y>�1� ?�)� �E{a�eЕ7D��1	�K��������y�v�Pb��;"ʪ7�� =��
#�ISs���`�7y�����:BsĢ�����sWM�-�4��YCZ����� u��&�#T���)�WꃭG�J���>������*x34}ζ��9쵥����$R /��%p�B�	y�V�I���PU\���C����4PVPm��5��L0�j"v��#/�>0�VI���
m���QG�;Y���}{�r����]�փ�oq���,*m����}����������a���4O��T����Q�Kl^�	&�l[
��Q�r�˨].�3�����j"i�7s��6x��.{�4᧊-��fKN-��e6��!���v��%�Q�hu"쒒�,�-*qH���o�����c:ӹb�S��� �����0��CSy���E��|���|@�����d
rG����[��k�l��K	�%�;��6'�V�U���[�V��k��n�!���V*BG���1�c|�Q.�X;k�͸�y�я�{c�������e���6X]	&ڀr�y��p�Ӂ��0� >�`w8��R�R|ؾ=��Ȉ���:��P����{��ƈ��}�Nƿ�|i�5��利ߑ��gD֔l��]��l�B�����|�y(�ǟ��7-�� z����J�1͠�]
�J��"f"8�O��*����t��m.*y$�%.w@a�W�B�:H-}��ԣyvr��F��8���Q1��ޖS�VO��QU�&���1-efSzC��~�~�=�����]S��Ky��_�����Z��u�g�dn�
Ji4�kyn�KW^+��h&���2'��|�2�$V�N"��^�?����;#�� !�aV��g�F���
zr�y<U�I@�Г��g��E�CR/
1~�<�ʨw��pp':SӴ��ǯ��쪏K58�_�0n���K"�!�^���{�����n�� ��@tK��h�p/=�9���k-OI�����]n
ܞW��I`�|�r���E�/櫪�V���,�X�b��w�w�7�_�l��g�6��h%Q���3��+�t�h�_�CH�Ì�j��8�/�Ѽ�{?�Ju�:�'v����Q�J�}���/[�	~cԈ��Pv>\�c����C��3�$����"�]���m��o[[��&��4�+��j%�)T��+��b^#;-�cr�c��Ϟ�"��wIi��x�,��m�\0_��1냥�Y9S�j�I��̴'���9m4/4��_���u��	!���/g��g�C�>�m<�K��B���*rN_J�۝fH��V�D�^�8J�s� ����2�>/FC;�&�O��'5��������r�퉛��7��@1��z�<�m�BAf���`��_18jR݀VCi�*㏨�x��a�g~M6���tS���v�J��]�ꭢ+2���pA�/Iw���I}u<�ƾ΄�_�dx���C[\��5,�8ܙ�6����2S�6��;җ���w>r��� ��|g�i